module SIMON_enc ( 
Kin_0,
Kin_1,
Kin_2,
Kin_3,
Kin_4,
Kin_5,
Kin_6,
Kin_7,
Kin_8,
Kin_9,
Kin_10,
Kin_11,
Kin_12,
Kin_13,
Kin_14,
Kin_15,
Kin_16,
Kin_17,
Kin_18,
Kin_19,
Kin_20,
Kin_21,
Kin_22,
Kin_23,
Kin_24,
Kin_25,
Kin_26,
Kin_27,
Kin_28,
Kin_29,
Kin_30,
Kin_31,
Kin_32,
Kin_33,
Kin_34,
Kin_35,
Kin_36,
Kin_37,
Kin_38,
Kin_39,
Kin_40,
Kin_41,
Kin_42,
Kin_43,
Kin_44,
Kin_45,
Kin_46,
Kin_47,
Kin_48,
Kin_49,
Kin_50,
Kin_51,
Kin_52,
Kin_53,
Kin_54,
Kin_55,
Kin_56,
Kin_57,
Kin_58,
Kin_59,
Kin_60,
Kin_61,
Kin_62,
Kin_63, 
Din_0,
Din_1,
Din_2,
Din_3,
Din_4,
Din_5,
Din_6,
Din_7,
Din_8,
Din_9,
Din_10,
Din_11,
Din_12,
Din_13,
Din_14,
Din_15,
Din_16,
Din_17,
Din_18,
Din_19,
Din_20,
Din_21,
Din_22,
Din_23,
Din_24,
Din_25,
Din_26,
Din_27,
Din_28,
Din_29,
Din_30,
Din_31,
Dout_0,
Dout_1,
Dout_2,
Dout_3,
Dout_4,
Dout_5,
Dout_6,
Dout_7,
Dout_8,
Dout_9,
Dout_10,
Dout_11,
Dout_12,
Dout_13,
Dout_14,
Dout_15,
Dout_16,
Dout_17,
Dout_18,
Dout_19,
Dout_20,
Dout_21,
Dout_22,
Dout_23,
Dout_24,
Dout_25,
Dout_26,
Dout_27,
Dout_28,
Dout_29,
Dout_30,
Dout_31,
Krdy, 
Drdy, 
Kvld, 
Dvld, 
EN, 
BSY, 
CLK, 
RSTn
);
//Start PIs
input Kin_0;
input Kin_1;
input Kin_2;
input Kin_3;
input Kin_4;
input Kin_5;
input Kin_6;
input Kin_7;
input Kin_8;
input Kin_9;
input Kin_10;
input Kin_11;
input Kin_12;
input Kin_13;
input Kin_14;
input Kin_15;
input Kin_16;
input Kin_17;
input Kin_18;
input Kin_19;
input Kin_20;
input Kin_21;
input Kin_22;
input Kin_23;
input Kin_24;
input Kin_25;
input Kin_26;
input Kin_27;
input Kin_28;
input Kin_29;
input Kin_30;
input Kin_31;
input Kin_32;
input Kin_33;
input Kin_34;
input Kin_35;
input Kin_36;
input Kin_37;
input Kin_38;
input Kin_39;
input Kin_40;
input Kin_41;
input Kin_42;
input Kin_43;
input Kin_44;
input Kin_45;
input Kin_46;
input Kin_47;
input Kin_48;
input Kin_49;
input Kin_50;
input Kin_51;
input Kin_52;
input Kin_53;
input Kin_54;
input Kin_55;
input Kin_56;
input Kin_57;
input Kin_58;
input Kin_59;
input Kin_60;
input Kin_61;
input Kin_62;
input Kin_63;
input Din_0;
input Din_1;
input Din_2;
input Din_3;
input Din_4;
input Din_5;
input Din_6;
input Din_7;
input Din_8;
input Din_9;
input Din_10;
input Din_11;
input Din_12;
input Din_13;
input Din_14;
input Din_15;
input Din_16;
input Din_17;
input Din_18;
input Din_19;
input Din_20;
input Din_21;
input Din_22;
input Din_23;
input Din_24;
input Din_25;
input Din_26;
input Din_27;
input Din_28;
input Din_29;
input Din_30;
input Din_31;
input Krdy;
input Drdy;
input EN; 
input CLK;
input RSTn;
//Start POs 
output Dout_0;
output Dout_1;
output Dout_2;
output Dout_3;
output Dout_4;
output Dout_5;
output Dout_6;
output Dout_7;
output Dout_8;
output Dout_9;
output Dout_10;
output Dout_11;
output Dout_12;
output Dout_13;
output Dout_14;
output Dout_15;
output Dout_16;
output Dout_17;
output Dout_18;
output Dout_19;
output Dout_20;
output Dout_21;
output Dout_22;
output Dout_23;
output Dout_24;
output Dout_25;
output Dout_26;
output Dout_27;
output Dout_28;
output Dout_29;
output Dout_30;
output Dout_31;
output Kvld;
output Dvld;
output BSY;
//Start wires
wire sel;
wire _keyexpantion_N27;
wire _keyexpantion_N26;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire rnd_0;
wire rnd_1;
wire rnd_2;
wire rnd_3;
wire rnd_4;
wire rnd_5;
wire rnd_6;
wire rnd_7;
wire rnd_8;
wire rnd_9;
wire rnd_10;
wire rnd_11;
wire rnd_12;
wire rnd_13;
wire rnd_14;
wire rnd_15;
wire rnd_16;
wire rnd_17;
wire rnd_18;
wire rnd_19;
wire rnd_20;
wire rnd_21;
wire rnd_22;
wire rnd_23;
wire rnd_24;
wire rnd_25;
wire rnd_26;
wire rnd_27;
wire rnd_28;
wire rnd_29;
wire rnd_30;
wire rnd_31;
wire dat_next_0;
wire dat_next_1;
wire dat_next_2;
wire dat_next_3;
wire dat_next_4;
wire dat_next_5;
wire dat_next_6;
wire dat_next_7;
wire dat_next_8;
wire dat_next_9;
wire dat_next_10;
wire dat_next_11;
wire dat_next_12;
wire dat_next_13;
wire dat_next_14;
wire dat_next_15;
wire dat_next_16;
wire dat_next_17;
wire dat_next_18;
wire dat_next_19;
wire dat_next_20;
wire dat_next_21;
wire dat_next_22;
wire dat_next_23;
wire dat_next_24;
wire dat_next_25;
wire dat_next_26;
wire dat_next_27;
wire dat_next_28;
wire dat_next_29;
wire dat_next_30;
wire dat_next_31;
wire rkey_next_0;
wire rkey_next_1;
wire rkey_next_2;
wire rkey_next_3;
wire rkey_next_4;
wire rkey_next_5;
wire rkey_next_6;
wire rkey_next_7;
wire rkey_next_8;
wire rkey_next_9;
wire rkey_next_10;
wire rkey_next_11;
wire rkey_next_12;
wire rkey_next_13;
wire rkey_next_14;
wire rkey_next_15;
wire rkey_next_16;
wire rkey_next_17;
wire rkey_next_18;
wire rkey_next_19;
wire rkey_next_20;
wire rkey_next_21;
wire rkey_next_22;
wire rkey_next_23;
wire rkey_next_24;
wire rkey_next_25;
wire rkey_next_26;
wire rkey_next_27;
wire rkey_next_28;
wire rkey_next_29;
wire rkey_next_30;
wire rkey_next_31;
wire rkey_next_32;
wire rkey_next_33;
wire rkey_next_34;
wire rkey_next_35;
wire rkey_next_36;
wire rkey_next_37;
wire rkey_next_38;
wire rkey_next_39;
wire rkey_next_40;
wire rkey_next_41;
wire rkey_next_42;
wire rkey_next_43;
wire rkey_next_44;
wire rkey_next_45;
wire rkey_next_46;
wire rkey_next_47;
wire rkey_next_48;
wire rkey_next_49;
wire rkey_next_50;
wire rkey_next_51;
wire rkey_next_52;
wire rkey_next_53;
wire rkey_next_54;
wire rkey_next_55;
wire rkey_next_56;
wire rkey_next_57;
wire rkey_next_58;
wire rkey_next_59;
wire rkey_next_60;
wire rkey_next_61;
wire rkey_next_62;
wire rkey_next_63;
wire rkey_0;
wire rkey_1;
wire rkey_2;
wire rkey_3;
wire rkey_4;
wire rkey_5;
wire rkey_6;
wire rkey_7;
wire rkey_8;
wire rkey_9;
wire rkey_10;
wire rkey_11;
wire rkey_12;
wire rkey_13;
wire rkey_14;
wire rkey_15;
wire rkey_16;
wire rkey_17;
wire rkey_18;
wire rkey_19;
wire rkey_20;
wire rkey_21;
wire rkey_22;
wire rkey_23;
wire rkey_24;
wire rkey_25;
wire rkey_26;
wire rkey_27;
wire rkey_28;
wire rkey_29;
wire rkey_30;
wire rkey_31;
wire rkey_32;
wire rkey_33;
wire rkey_34;
wire rkey_35;
wire rkey_36;
wire rkey_37;
wire rkey_38;
wire rkey_39;
wire rkey_40;
wire rkey_41;
wire rkey_42;
wire rkey_43;
wire rkey_44;
wire rkey_45;
wire rkey_46;
wire rkey_47;
wire rkey_48;
wire rkey_49;
wire rkey_50;
wire rkey_51;
wire rkey_52;
wire rkey_53;
wire rkey_54;
wire rkey_55;
wire rkey_56;
wire rkey_57;
wire rkey_58;
wire rkey_59;
wire rkey_60;
wire rkey_61;
wire rkey_62;
wire rkey_63;
wire key_0;
wire key_1;
wire key_2;
wire key_3;
wire key_4;
wire key_5;
wire key_6;
wire key_7;
wire key_8;
wire key_9;
wire key_10;
wire key_11;
wire key_12;
wire key_13;
wire key_14;
wire key_15;
wire key_16;
wire key_17;
wire key_18;
wire key_19;
wire key_20;
wire key_21;
wire key_22;
wire key_23;
wire key_24;
wire key_25;
wire key_26;
wire key_27;
wire key_28;
wire key_29;
wire key_30;
wire key_31;
wire key_32;
wire key_33;
wire key_34;
wire key_35;
wire key_36;
wire key_37;
wire key_38;
wire key_39;
wire key_40;
wire key_41;
wire key_42;
wire key_43;
wire key_44;
wire key_45;
wire key_46;
wire key_47;
wire key_48;
wire key_49;
wire key_50;
wire key_51;
wire key_52;
wire key_53;
wire key_54;
wire key_55;
wire key_56;
wire key_57;
wire key_58;
wire key_59;
wire key_60;
wire key_61;
wire key_62;
wire key_63;
//Start cells
  QDFFRBHHD Kvld_reg ( .D(n483), .CK(CLK), .RB(RSTn), .Q(Kvld) );
  QDFFRBHHD sel_reg ( .D(n482), .CK(CLK), .RB(RSTn), .Q(sel) );
  QDFFRBHHD Dvld_reg ( .D(n481), .CK(CLK), .RB(RSTn), .Q(Dvld) );
  QDFFRBHHD BSY_reg ( .D(n480), .CK(CLK), .RB(RSTn), .Q(BSY) );
  QDFFRBHHD _rkey_reg_0  ( .D(n479), .CK(CLK), .RB(RSTn), .Q(rkey_0) );
  QDFFRBHHD _rkey_reg_48  ( .D(n478), .CK(CLK), .RB(RSTn), .Q(rkey_next_32));
  QDFFRBHHD _rkey_reg_32  ( .D(n477), .CK(CLK), .RB(RSTn), .Q(rkey_next_16));
  QDFFRBHHD _rkey_reg_16  ( .D(n476), .CK(CLK), .RB(RSTn), .Q(rkey_next_0));
  QDFFRBHHD _rkey_reg_61  ( .D(n475), .CK(CLK), .RB(RSTn), .Q(rkey_next_45));
  QDFFRBHHD _rkey_reg_45  ( .D(n474), .CK(CLK), .RB(RSTn), .Q(rkey_next_29));
  QDFFRBHHD _rkey_reg_29  ( .D(n473), .CK(CLK), .RB(RSTn), .Q(rkey_next_13));
  QDFFRBHHD _rkey_reg_13  ( .D(n472), .CK(CLK), .RB(RSTn), .Q(rkey_13) );
  QDFFRBHHD _rkey_reg_58  ( .D(n471), .CK(CLK), .RB(RSTn), .Q(rkey_next_42));
  QDFFRBHHD _rkey_reg_42  ( .D(n470), .CK(CLK), .RB(RSTn), .Q(rkey_next_26));
  QDFFRBHHD _rkey_reg_26  ( .D(n469), .CK(CLK), .RB(RSTn), .Q(rkey_next_10));
  QDFFRBHHD _rkey_reg_10  ( .D(n468), .CK(CLK), .RB(RSTn), .Q(rkey_10) );
  QDFFRBHHD _rkey_reg_55  ( .D(n467), .CK(CLK), .RB(RSTn), .Q(rkey_next_39));
  QDFFRBHHD _rkey_reg_39  ( .D(n466), .CK(CLK), .RB(RSTn), .Q(rkey_next_23));
  QDFFRBHHD _rkey_reg_23  ( .D(n465), .CK(CLK), .RB(RSTn), .Q(rkey_next_7));
  QDFFRBHHD _rkey_reg_7  ( .D(n464), .CK(CLK), .RB(RSTn), .Q(rkey_7) );
  QDFFRBHHD _rkey_reg_52  ( .D(n463), .CK(CLK), .RB(RSTn), .Q(rkey_next_36));
  QDFFRBHHD _rkey_reg_36  ( .D(n462), .CK(CLK), .RB(RSTn), .Q(rkey_next_20));
  QDFFRBHHD _rkey_reg_20  ( .D(n461), .CK(CLK), .RB(RSTn), .Q(rkey_next_4));
  QDFFRBHHD _rkey_reg_4  ( .D(n460), .CK(CLK), .RB(RSTn), .Q(rkey_4) );
  QDFFRBHHD _rkey_reg_49  ( .D(n459), .CK(CLK), .RB(RSTn), .Q(rkey_next_33));
  QDFFRBHHD _rkey_reg_33  ( .D(n458), .CK(CLK), .RB(RSTn), .Q(rkey_next_17));
  QDFFRBHHD _rkey_reg_17  ( .D(n457), .CK(CLK), .RB(RSTn), .Q(rkey_next_1));
  QDFFRBHHD _rkey_reg_1  ( .D(n456), .CK(CLK), .RB(RSTn), .Q(rkey_1) );
  QDFFRBHHD _rkey_reg_62  ( .D(n455), .CK(CLK), .RB(RSTn), .Q(rkey_next_46));
  QDFFRBHHD _rkey_reg_46  ( .D(n454), .CK(CLK), .RB(RSTn), .Q(rkey_next_30));
  QDFFRBHHD _rkey_reg_30  ( .D(n453), .CK(CLK), .RB(RSTn), .Q(rkey_next_14));
  QDFFRBHHD _rkey_reg_14  ( .D(n452), .CK(CLK), .RB(RSTn), .Q(rkey_14) );
  QDFFRBHHD _rkey_reg_59  ( .D(n451), .CK(CLK), .RB(RSTn), .Q(rkey_next_43));
  QDFFRBHHD _rkey_reg_43  ( .D(n450), .CK(CLK), .RB(RSTn), .Q(rkey_next_27));
  QDFFRBHHD _rkey_reg_27  ( .D(n449), .CK(CLK), .RB(RSTn), .Q(rkey_next_11));
  QDFFRBHHD _rkey_reg_11  ( .D(n448), .CK(CLK), .RB(RSTn), .Q(rkey_11) );
  QDFFRBHHD _rkey_reg_56  ( .D(n447), .CK(CLK), .RB(RSTn), .Q(rkey_next_40));
  QDFFRBHHD _rkey_reg_40  ( .D(n446), .CK(CLK), .RB(RSTn), .Q(rkey_next_24));
  QDFFRBHHD _rkey_reg_24  ( .D(n445), .CK(CLK), .RB(RSTn), .Q(rkey_next_8));
  QDFFRBHHD _rkey_reg_8  ( .D(n444), .CK(CLK), .RB(RSTn), .Q(rkey_8) );
  QDFFRBHHD _rkey_reg_53  ( .D(n443), .CK(CLK), .RB(RSTn), .Q(rkey_next_37));
  QDFFRBHHD _rkey_reg_37  ( .D(n442), .CK(CLK), .RB(RSTn), .Q(rkey_next_21));
  QDFFRBHHD _rkey_reg_21  ( .D(n441), .CK(CLK), .RB(RSTn), .Q(rkey_next_5));
  QDFFRBHHD _rkey_reg_5  ( .D(n440), .CK(CLK), .RB(RSTn), .Q(rkey_5) );
  QDFFRBHHD _rkey_reg_50  ( .D(n439), .CK(CLK), .RB(RSTn), .Q(rkey_next_34));
  QDFFRBHHD _rkey_reg_34  ( .D(n438), .CK(CLK), .RB(RSTn), .Q(rkey_next_18));
  QDFFRBHHD _rkey_reg_18  ( .D(n437), .CK(CLK), .RB(RSTn), .Q(rkey_next_2));
  QDFFRBHHD _rkey_reg_2  ( .D(n436), .CK(CLK), .RB(RSTn), .Q(rkey_2) );
  QDFFRBHHD _rkey_reg_63  ( .D(n435), .CK(CLK), .RB(RSTn), .Q(rkey_next_47));
  QDFFRBHHD _rkey_reg_47  ( .D(n434), .CK(CLK), .RB(RSTn), .Q(rkey_next_31));
  QDFFRBHHD _rkey_reg_31  ( .D(n433), .CK(CLK), .RB(RSTn), .Q(rkey_next_15));
  QDFFRBHHD _rkey_reg_15  ( .D(n432), .CK(CLK), .RB(RSTn), .Q(rkey_15) );
  QDFFRBHHD _rkey_reg_60  ( .D(n431), .CK(CLK), .RB(RSTn), .Q(rkey_next_44));
  QDFFRBHHD _rkey_reg_44  ( .D(n430), .CK(CLK), .RB(RSTn), .Q(rkey_next_28));
  QDFFRBHHD _rkey_reg_28  ( .D(n429), .CK(CLK), .RB(RSTn), .Q(rkey_next_12));
  QDFFRBHHD _rkey_reg_12  ( .D(n428), .CK(CLK), .RB(RSTn), .Q(rkey_12) );
  QDFFRBHHD _rkey_reg_57  ( .D(n427), .CK(CLK), .RB(RSTn), .Q(rkey_next_41));
  QDFFRBHHD _rkey_reg_41  ( .D(n426), .CK(CLK), .RB(RSTn), .Q(rkey_next_25));
  QDFFRBHHD _rkey_reg_25  ( .D(n425), .CK(CLK), .RB(RSTn), .Q(rkey_next_9));
  QDFFRBHHD _rkey_reg_9  ( .D(n424), .CK(CLK), .RB(RSTn), .Q(rkey_9) );
  QDFFRBHHD _rkey_reg_54  ( .D(n423), .CK(CLK), .RB(RSTn), .Q(rkey_next_38));
  QDFFRBHHD _rkey_reg_38  ( .D(n422), .CK(CLK), .RB(RSTn), .Q(rkey_next_22));
  QDFFRBHHD _rkey_reg_22  ( .D(n421), .CK(CLK), .RB(RSTn), .Q(rkey_next_6));
  QDFFRBHHD _rkey_reg_6  ( .D(n420), .CK(CLK), .RB(RSTn), .Q(rkey_6) );
  QDFFRBHHD _rkey_reg_51  ( .D(n419), .CK(CLK), .RB(RSTn), .Q(rkey_next_35));
  QDFFRBHHD _rkey_reg_35  ( .D(n418), .CK(CLK), .RB(RSTn), .Q(rkey_next_19));
  QDFFRBHHD _rkey_reg_19  ( .D(n417), .CK(CLK), .RB(RSTn), .Q(rkey_next_3));
  QDFFRBHHD _rkey_reg_3  ( .D(n416), .CK(CLK), .RB(RSTn), .Q(rkey_3) );
  QDFFRBHHD _rnd_reg_1  ( .D(n610), .CK(CLK), .RB(RSTn), .Q(_keyexpantion_N27 ) );
  QDFFRBHHD _rnd_reg_2  ( .D(n609), .CK(CLK), .RB(RSTn), .Q(rnd_2) );
  QDFFRBHHD _rnd_reg_3  ( .D(n608), .CK(CLK), .RB(RSTn), .Q(rnd_3) );
  QDFFRBHHD _rnd_reg_4  ( .D(n607), .CK(CLK), .RB(RSTn), .Q(rnd_4) );
  QDFFRBHHD _rnd_reg_5  ( .D(n606), .CK(CLK), .RB(RSTn), .Q(rnd_5) );
  QDFFRBHHD _rnd_reg_6  ( .D(n605), .CK(CLK), .RB(RSTn), .Q(rnd_6) );
  QDFFRBHHD _rnd_reg_7  ( .D(n604), .CK(CLK), .RB(RSTn), .Q(rnd_7) );
  QDFFRBHHD _rnd_reg_8  ( .D(n603), .CK(CLK), .RB(RSTn), .Q(rnd_8) );
  QDFFRBHHD _rnd_reg_9  ( .D(n602), .CK(CLK), .RB(RSTn), .Q(rnd_9) );
  QDFFRBHHD _rnd_reg_10  ( .D(n601), .CK(CLK), .RB(RSTn), .Q(rnd_10) );
  QDFFRBHHD _rnd_reg_11  ( .D(n600), .CK(CLK), .RB(RSTn), .Q(rnd_11) );
  QDFFRBHHD _rnd_reg_12  ( .D(n599), .CK(CLK), .RB(RSTn), .Q(rnd_12) );
  QDFFRBHHD _rnd_reg_13  ( .D(n598), .CK(CLK), .RB(RSTn), .Q(rnd_13) );
  QDFFRBHHD _rnd_reg_14  ( .D(n597), .CK(CLK), .RB(RSTn), .Q(rnd_14) );
  QDFFRBHHD _rnd_reg_15  ( .D(n596), .CK(CLK), .RB(RSTn), .Q(rnd_15) );
  QDFFRBHHD _rnd_reg_16  ( .D(n595), .CK(CLK), .RB(RSTn), .Q(rnd_16) );
  QDFFRBHHD _rnd_reg_17  ( .D(n594), .CK(CLK), .RB(RSTn), .Q(rnd_17) );
  QDFFRBHHD _rnd_reg_18  ( .D(n593), .CK(CLK), .RB(RSTn), .Q(rnd_18) );
  QDFFRBHHD _rnd_reg_19  ( .D(n592), .CK(CLK), .RB(RSTn), .Q(rnd_19) );
  QDFFRBHHD _rnd_reg_20  ( .D(n591), .CK(CLK), .RB(RSTn), .Q(rnd_20) );
  QDFFRBHHD _rnd_reg_21  ( .D(n590), .CK(CLK), .RB(RSTn), .Q(rnd_21) );
  QDFFRBHHD _rnd_reg_22  ( .D(n589), .CK(CLK), .RB(RSTn), .Q(rnd_22) );
  QDFFRBHHD _rnd_reg_23  ( .D(n588), .CK(CLK), .RB(RSTn), .Q(rnd_23) );
  QDFFRBHHD _rnd_reg_24  ( .D(n587), .CK(CLK), .RB(RSTn), .Q(rnd_24) );
  QDFFRBHHD _rnd_reg_25  ( .D(n586), .CK(CLK), .RB(RSTn), .Q(rnd_25) );
  QDFFRBHHD _rnd_reg_26  ( .D(n585), .CK(CLK), .RB(RSTn), .Q(rnd_26) );
  QDFFRBHHD _rnd_reg_27  ( .D(n584), .CK(CLK), .RB(RSTn), .Q(rnd_27) );
  QDFFRBHHD _rnd_reg_28  ( .D(n583), .CK(CLK), .RB(RSTn), .Q(rnd_28) );
  QDFFRBHHD _rnd_reg_29  ( .D(n582), .CK(CLK), .RB(RSTn), .Q(rnd_29) );
  QDFFRBHHD _rnd_reg_30  ( .D(n581), .CK(CLK), .RB(RSTn), .Q(rnd_30) );
  QDFFRBHHD _rnd_reg_31  ( .D(n612), .CK(CLK), .RB(RSTn), .Q(rnd_31) );
  QDFFRBHHD _key_reg_63  ( .D(n580), .CK(CLK), .RB(RSTn), .Q(key_63) );
  QDFFRBHHD _key_reg_62  ( .D(n579), .CK(CLK), .RB(RSTn), .Q(key_62) );
  QDFFRBHHD _key_reg_61  ( .D(n578), .CK(CLK), .RB(RSTn), .Q(key_61) );
  QDFFRBHHD _key_reg_60  ( .D(n577), .CK(CLK), .RB(RSTn), .Q(key_60) );
  QDFFRBHHD _key_reg_59  ( .D(n576), .CK(CLK), .RB(RSTn), .Q(key_59) );
  QDFFRBHHD _key_reg_58  ( .D(n575), .CK(CLK), .RB(RSTn), .Q(key_58) );
  QDFFRBHHD _key_reg_57  ( .D(n574), .CK(CLK), .RB(RSTn), .Q(key_57) );
  QDFFRBHHD _key_reg_56  ( .D(n573), .CK(CLK), .RB(RSTn), .Q(key_56) );
  QDFFRBHHD _key_reg_55  ( .D(n572), .CK(CLK), .RB(RSTn), .Q(key_55) );
  QDFFRBHHD _key_reg_54  ( .D(n571), .CK(CLK), .RB(RSTn), .Q(key_54) );
  QDFFRBHHD _key_reg_53  ( .D(n570), .CK(CLK), .RB(RSTn), .Q(key_53) );
  QDFFRBHHD _key_reg_52  ( .D(n569), .CK(CLK), .RB(RSTn), .Q(key_52) );
  QDFFRBHHD _key_reg_51  ( .D(n568), .CK(CLK), .RB(RSTn), .Q(key_51) );
  QDFFRBHHD _key_reg_50  ( .D(n567), .CK(CLK), .RB(RSTn), .Q(key_50) );
  QDFFRBHHD _key_reg_49  ( .D(n566), .CK(CLK), .RB(RSTn), .Q(key_49) );
  QDFFRBHHD _key_reg_48  ( .D(n565), .CK(CLK), .RB(RSTn), .Q(key_48) );
  QDFFRBHHD _key_reg_47  ( .D(n564), .CK(CLK), .RB(RSTn), .Q(key_47) );
  QDFFRBHHD _key_reg_46  ( .D(n563), .CK(CLK), .RB(RSTn), .Q(key_46) );
  QDFFRBHHD _key_reg_45  ( .D(n562), .CK(CLK), .RB(RSTn), .Q(key_45) );
  QDFFRBHHD _key_reg_44  ( .D(n561), .CK(CLK), .RB(RSTn), .Q(key_44) );
  QDFFRBHHD _key_reg_43  ( .D(n560), .CK(CLK), .RB(RSTn), .Q(key_43) );
  QDFFRBHHD _key_reg_42  ( .D(n559), .CK(CLK), .RB(RSTn), .Q(key_42) );
  QDFFRBHHD _key_reg_41  ( .D(n558), .CK(CLK), .RB(RSTn), .Q(key_41) );
  QDFFRBHHD _key_reg_40  ( .D(n557), .CK(CLK), .RB(RSTn), .Q(key_40) );
  QDFFRBHHD _key_reg_39  ( .D(n556), .CK(CLK), .RB(RSTn), .Q(key_39) );
  QDFFRBHHD _key_reg_38  ( .D(n555), .CK(CLK), .RB(RSTn), .Q(key_38) );
  QDFFRBHHD _key_reg_37  ( .D(n554), .CK(CLK), .RB(RSTn), .Q(key_37) );
  QDFFRBHHD _key_reg_36  ( .D(n553), .CK(CLK), .RB(RSTn), .Q(key_36) );
  QDFFRBHHD _key_reg_35  ( .D(n552), .CK(CLK), .RB(RSTn), .Q(key_35) );
  QDFFRBHHD _key_reg_34  ( .D(n551), .CK(CLK), .RB(RSTn), .Q(key_34) );
  QDFFRBHHD _key_reg_33  ( .D(n550), .CK(CLK), .RB(RSTn), .Q(key_33) );
  QDFFRBHHD _key_reg_32  ( .D(n549), .CK(CLK), .RB(RSTn), .Q(key_32) );
  QDFFRBHHD _key_reg_31  ( .D(n548), .CK(CLK), .RB(RSTn), .Q(key_31) );
  QDFFRBHHD _key_reg_30  ( .D(n547), .CK(CLK), .RB(RSTn), .Q(key_30) );
  QDFFRBHHD _key_reg_29  ( .D(n546), .CK(CLK), .RB(RSTn), .Q(key_29) );
  QDFFRBHHD _key_reg_28  ( .D(n545), .CK(CLK), .RB(RSTn), .Q(key_28) );
  QDFFRBHHD _key_reg_27  ( .D(n544), .CK(CLK), .RB(RSTn), .Q(key_27) );
  QDFFRBHHD _key_reg_26  ( .D(n543), .CK(CLK), .RB(RSTn), .Q(key_26) );
  QDFFRBHHD _key_reg_25  ( .D(n542), .CK(CLK), .RB(RSTn), .Q(key_25) );
  QDFFRBHHD _key_reg_24  ( .D(n541), .CK(CLK), .RB(RSTn), .Q(key_24) );
  QDFFRBHHD _key_reg_23  ( .D(n540), .CK(CLK), .RB(RSTn), .Q(key_23) );
  QDFFRBHHD _key_reg_22  ( .D(n539), .CK(CLK), .RB(RSTn), .Q(key_22) );
  QDFFRBHHD _key_reg_21  ( .D(n538), .CK(CLK), .RB(RSTn), .Q(key_21) );
  QDFFRBHHD _key_reg_20  ( .D(n537), .CK(CLK), .RB(RSTn), .Q(key_20) );
  QDFFRBHHD _key_reg_19  ( .D(n536), .CK(CLK), .RB(RSTn), .Q(key_19) );
  QDFFRBHHD _key_reg_18  ( .D(n535), .CK(CLK), .RB(RSTn), .Q(key_18) );
  QDFFRBHHD _key_reg_17  ( .D(n534), .CK(CLK), .RB(RSTn), .Q(key_17) );
  QDFFRBHHD _key_reg_16  ( .D(n533), .CK(CLK), .RB(RSTn), .Q(key_16) );
  QDFFRBHHD _key_reg_15  ( .D(n532), .CK(CLK), .RB(RSTn), .Q(key_15) );
  QDFFRBHHD _key_reg_14  ( .D(n531), .CK(CLK), .RB(RSTn), .Q(key_14) );
  QDFFRBHHD _key_reg_13  ( .D(n530), .CK(CLK), .RB(RSTn), .Q(key_13) );
  QDFFRBHHD _key_reg_12  ( .D(n529), .CK(CLK), .RB(RSTn), .Q(key_12) );
  QDFFRBHHD _key_reg_11  ( .D(n528), .CK(CLK), .RB(RSTn), .Q(key_11) );
  QDFFRBHHD _key_reg_10  ( .D(n527), .CK(CLK), .RB(RSTn), .Q(key_10) );
  QDFFRBHHD _key_reg_9  ( .D(n526), .CK(CLK), .RB(RSTn), .Q(key_9) );
  QDFFRBHHD _key_reg_8  ( .D(n525), .CK(CLK), .RB(RSTn), .Q(key_8) );
  QDFFRBHHD _key_reg_7  ( .D(n524), .CK(CLK), .RB(RSTn), .Q(key_7) );
  QDFFRBHHD _key_reg_6  ( .D(n523), .CK(CLK), .RB(RSTn), .Q(key_6) );
  QDFFRBHHD _key_reg_5  ( .D(n522), .CK(CLK), .RB(RSTn), .Q(key_5) );
  QDFFRBHHD _key_reg_4  ( .D(n521), .CK(CLK), .RB(RSTn), .Q(key_4) );
  QDFFRBHHD _key_reg_3  ( .D(n520), .CK(CLK), .RB(RSTn), .Q(key_3) );
  QDFFRBHHD _key_reg_2  ( .D(n519), .CK(CLK), .RB(RSTn), .Q(key_2) );
  QDFFRBHHD _key_reg_1  ( .D(n518), .CK(CLK), .RB(RSTn), .Q(key_1) );
  QDFFRBHHD _key_reg_0  ( .D(n517), .CK(CLK), .RB(RSTn), .Q(key_0) );
  QDFFRBHHD _dat_reg_16  ( .D(n500), .CK(CLK), .RB(RSTn), .Q(dat_next_0) );
  QDFFRBHHD _dat_reg_0  ( .D(n516), .CK(CLK), .RB(RSTn), .Q(Dout_0) );
  QDFFRBHHD _dat_reg_24  ( .D(n492), .CK(CLK), .RB(RSTn), .Q(dat_next_8) );
  QDFFRBHHD _dat_reg_8  ( .D(n508), .CK(CLK), .RB(RSTn), .Q(Dout_8) );
  QDFFRBHHD _dat_reg_26  ( .D(n490), .CK(CLK), .RB(RSTn), .Q(dat_next_10) );
  QDFFRBHHD _dat_reg_10  ( .D(n506), .CK(CLK), .RB(RSTn), .Q(Dout_10) );
  QDFFRBHHD _dat_reg_28  ( .D(n488), .CK(CLK), .RB(RSTn), .Q(dat_next_12) );
  QDFFRBHHD _dat_reg_12  ( .D(n504), .CK(CLK), .RB(RSTn), .Q(Dout_12) );
  QDFFRBHHD _dat_reg_30  ( .D(n486), .CK(CLK), .RB(RSTn), .Q(dat_next_14) );
  QDFFRBHHD _dat_reg_14  ( .D(n502), .CK(CLK), .RB(RSTn), .Q(Dout_14) );
  QDFFRBHHD _dat_reg_31  ( .D(n484), .CK(CLK), .RB(RSTn), .Q(dat_next_15) );
  QDFFRBHHD _dat_reg_15  ( .D(n501), .CK(CLK), .RB(RSTn), .Q(Dout_15) );
  QDFFRBHHD _dat_reg_23  ( .D(n493), .CK(CLK), .RB(RSTn), .Q(dat_next_7) );
  QDFFRBHHD _dat_reg_7  ( .D(n509), .CK(CLK), .RB(RSTn), .Q(Dout_7) );
  QDFFRBHHD _dat_reg_25  ( .D(n491), .CK(CLK), .RB(RSTn), .Q(dat_next_9) );
  QDFFRBHHD _dat_reg_9  ( .D(n507), .CK(CLK), .RB(RSTn), .Q(Dout_9) );
  QDFFRBHHD _dat_reg_17  ( .D(n499), .CK(CLK), .RB(RSTn), .Q(dat_next_1) );
  QDFFRBHHD _dat_reg_1  ( .D(n515), .CK(CLK), .RB(RSTn), .Q(Dout_1) );
  QDFFRBHHD _dat_reg_18  ( .D(n498), .CK(CLK), .RB(RSTn), .Q(dat_next_2) );
  QDFFRBHHD _dat_reg_2  ( .D(n514), .CK(CLK), .RB(RSTn), .Q(Dout_2) );
  QDFFRBHHD _dat_reg_27  ( .D(n489), .CK(CLK), .RB(RSTn), .Q(dat_next_11) );
  QDFFRBHHD _dat_reg_11  ( .D(n505), .CK(CLK), .RB(RSTn), .Q(Dout_11) );
  QDFFRBHHD _dat_reg_19  ( .D(n497), .CK(CLK), .RB(RSTn), .Q(dat_next_3) );
  QDFFRBHHD _dat_reg_3  ( .D(n513), .CK(CLK), .RB(RSTn), .Q(Dout_3) );
  QDFFRBHHD _dat_reg_20  ( .D(n496), .CK(CLK), .RB(RSTn), .Q(dat_next_4) );
  QDFFRBHHD _dat_reg_4  ( .D(n512), .CK(CLK), .RB(RSTn), .Q(Dout_4) );
  QDFFRBHHD _dat_reg_29  ( .D(n487), .CK(CLK), .RB(RSTn), .Q(dat_next_13) );
  QDFFRBHHD _dat_reg_13  ( .D(n503), .CK(CLK), .RB(RSTn), .Q(Dout_13) );
  QDFFRBHHD _dat_reg_21  ( .D(n495), .CK(CLK), .RB(RSTn), .Q(dat_next_5) );
  QDFFRBHHD _dat_reg_5  ( .D(n511), .CK(CLK), .RB(RSTn), .Q(Dout_5) );
  QDFFRBHHD _dat_reg_22  ( .D(n494), .CK(CLK), .RB(RSTn), .Q(dat_next_6) );
  QDFFRBHHD _dat_reg_6  ( .D(n510), .CK(CLK), .RB(RSTn), .Q(Dout_6) );
  DFFSBEHD _rnd_reg_0  ( .D(n611), .CK(CLK), .SB(RSTn), .Q(_keyexpantion_N26 ), .QB(n1857) );
  INVDHD U616 ( .I(EN), .O(n1584) );
  INVDHD U617 ( .I(n734), .O(n652) );
  NR2EHD U618 ( .I1(n735), .I2(n724), .O(n723) );
  INVDHD U619 ( .I(n1291), .O(n1289) );
  XNR2EHD U620 ( .I1(n1217), .I2(n1216), .O(n1236) );
  INVDHD U621 ( .I(n1021), .O(n1028) );
  XNR2EHD U622 ( .I1(n1098), .I2(n1100), .O(n627) );
  INVDHD U623 ( .I(n681), .O(n849) );
  INVDHD U624 ( .I(n1250), .O(n660) );
  XNR2HHD U625 ( .I1(n1069), .I2(n1202), .O(n1118) );
  ND2CHD U626 ( .I1(n1006), .I2(rnd_28), .O(n1009) );
  XOR2EHD U627 ( .I1(rnd_25), .I2(n1073), .O(n1072) );
  INVGHD U628 ( .I(n1005), .O(n1092) );
  XNR2HHD U629 ( .I1(n1091), .I2(n1005), .O(n1144) );
  NR2GHD U630 ( .I1(n987), .I2(n1062), .O(n1000) );
  INVHHD U631 ( .I(n898), .O(n1061) );
  INVDHD U632 ( .I(n982), .O(n755) );
  XNR2HHD U633 ( .I1(rnd_15), .I2(n694), .O(n1039) );
  ND2DHD U634 ( .I1(n749), .I2(n787), .O(n748) );
  INVGHD U635 ( .I(rnd_2), .O(n1579) );
  BUFCKIHD U636 ( .I(n975), .O(n632) );
  INVGHD U637 ( .I(rnd_19), .O(n1561) );
  INVGHD U638 ( .I(rnd_20), .O(n1562) );
  INVLHD U639 ( .I(rnd_14), .O(n1350) );
  XNR2EHD U640 ( .I1(n1108), .I2(n621), .O(n1132) );
  ND2HHD U641 ( .I1(n750), .I2(n748), .O(n1140) );
  XNR2HHD U642 ( .I1(rnd_29), .I2(n1113), .O(n1252) );
  BUFEHD U643 ( .I(n1330), .O(n1852) );
  ND2DHD U644 ( .I1(n1349), .I2(EN), .O(n1570) );
  INVKHD U645 ( .I(n868), .O(n917) );
  INVLHD U646 ( .I(n1034), .O(n768) );
  ND2HHD U647 ( .I1(n1201), .I2(n1200), .O(n1235) );
  ND2HHD U648 ( .I1(n1255), .I2(n1114), .O(n1065) );
  INVDHD U649 ( .I(n1150), .O(n1153) );
  NR2GHD U650 ( .I1(rnd_19), .I2(rnd_18), .O(n934) );
  NR2EHD U651 ( .I1(n1148), .I2(n780), .O(n779) );
  MAO222EHD U652 ( .A1(n1147), .B1(n1146), .C1(n1145), .O(n1148) );
  NR2BHD U653 ( .I1(n789), .I2(n869), .O(n786) );
  ND2HHD U654 ( .I1(n1104), .I2(n1103), .O(n1151) );
  INVCHD U655 ( .I(n1047), .O(n1048) );
  AN2HHD U656 ( .I1(n1074), .I2(n719), .O(n1047) );
  INVGHD U657 ( .I(n758), .O(n733) );
  ND2DHD U658 ( .I1(n1030), .I2(n1031), .O(n741) );
  INVCKGHD U659 ( .I(n632), .O(n1319) );
  INVCKGHD U660 ( .I(n1222), .O(n683) );
  ND2HHD U661 ( .I1(n904), .I2(n923), .O(n907) );
  NR2CHD U662 ( .I1(n918), .I2(n1315), .O(n919) );
  OA12EHD U663 ( .B1(n992), .B2(n996), .A1(n995), .O(n1111) );
  XNR2KHD U664 ( .I1(n1082), .I2(n1081), .O(n1087) );
  ND2HHD U665 ( .I1(n892), .I2(n891), .O(n906) );
  INVGHD U666 ( .I(n1163), .O(n614) );
  AOI22BHD U667 ( .A1(Din_16), .A2(n1573), .B1(n1571), .B2(dat_next_0), .O(n1299) );
  ND2DHD U668 ( .I1(n1298), .I2(EN), .O(n1571) );
  NR2CHD U669 ( .I1(n1577), .I2(n1578), .O(n1845) );
  NR2CHD U670 ( .I1(n1579), .I2(n1578), .O(n1851) );
  MXL2CHD U671 ( .A(n1561), .B(n1562), .S(n1570), .OB(n591) );
  MXL2CHD U672 ( .A(n1560), .B(n1561), .S(n1570), .OB(n592) );
  XNR2CHD U673 ( .I1(rnd_7), .I2(n746), .O(n745) );
  AN2HHD U674 ( .I1(n1297), .I2(n1295), .O(n1572) );
  ND2DHD U675 ( .I1(n1583), .I2(n1553), .O(n1578) );
  AN2EHD U676 ( .I1(_keyexpantion_N27 ), .I2(n1583), .O(n1844) );
  ND2DHD U677 ( .I1(n1294), .I2(_keyexpantion_N26 ), .O(n1297) );
  NR2CHD U678 ( .I1(n1328), .I2(_keyexpantion_N26 ), .O(n1583) );
  INVDHD U679 ( .I(_keyexpantion_N27 ), .O(n1553) );
  ND2DHD U680 ( .I1(_keyexpantion_N26 ), .I2(n1348), .O(n1349) );
  INVGHD U681 ( .I(rnd_6), .O(n914) );
  NR2CHD U682 ( .I1(Drdy), .I2(n1584), .O(n1295) );
  ND2DHD U683 ( .I1(n1327), .I2(EN), .O(n1328) );
  AN2EHD U684 ( .I1(EN), .I2(Drdy), .O(n1573) );
  AN2HHD U685 ( .I1(EN), .I2(Krdy), .O(n1807) );
  XNR2HHD U686 ( .I1(n1129), .I2(n1126), .O(n780) );
  OR2EHD U687 ( .I1(n1022), .I2(n785), .O(n617) );
  ND2HHD U688 ( .I1(n861), .I2(n860), .O(n862) );
  BUFLHD U689 ( .I(n975), .O(n878) );
  ND2HHD U690 ( .I1(n740), .I2(n991), .O(n998) );
  ND2HHD U691 ( .I1(n1115), .I2(n1202), .O(n848) );
  NR2IHD U692 ( .I1(rnd_14), .I2(n1115), .O(n681) );
  INVGHD U693 ( .I(n1115), .O(n1255) );
  INVCKGHD U694 ( .I(n965), .O(n966) );
  XNR2KHD U695 ( .I1(rnd_31), .I2(n876), .O(n896) );
  NR2GHD U696 ( .I1(_keyexpantion_N26 ), .I2(n1137), .O(n990) );
  INVGHD U697 ( .I(n1143), .O(n997) );
  INVCKGHD U698 ( .I(n1110), .O(n984) );
  NR2CHD U699 ( .I1(n1163), .I2(n758), .O(n757) );
  INVHHD U700 ( .I(n988), .O(n999) );
  INVHHD U701 ( .I(n842), .O(n1329) );
  NR2GHD U702 ( .I1(n852), .I2(n1034), .O(n877) );
  NR2GHD U703 ( .I1(n1033), .I2(n1034), .O(n821) );
  NR2GHD U704 ( .I1(rnd_18), .I2(n1034), .O(n794) );
  ND2HHD U705 ( .I1(n638), .I2(n637), .O(n959) );
  ND2DHD U706 ( .I1(n882), .I2(n881), .O(n886) );
  INVGHD U707 ( .I(n1114), .O(n1066) );
  NR2EHD U708 ( .I1(n875), .I2(n1034), .O(n876) );
  INVLHD U709 ( .I(n820), .O(n1034) );
  ND2DHD U710 ( .I1(n951), .I2(n997), .O(n955) );
  XNR2HHD U711 ( .I1(n1143), .I2(n698), .O(n1041) );
  NR2EHD U712 ( .I1(n910), .I2(n1034), .O(n773) );
  XNR2HHD U713 ( .I1(n1560), .I2(n1034), .O(n1005) );
  INVDHD U714 ( .I(n1270), .O(n1275) );
  AN2HHD U715 ( .I1(n1272), .I2(n1270), .O(n615) );
  ND2HHD U716 ( .I1(n658), .I2(n1183), .O(n642) );
  ND2DHD U717 ( .I1(n1239), .I2(n1566), .O(n861) );
  INVDHD U718 ( .I(n1215), .O(n1239) );
  ND3CHD U719 ( .I1(n766), .I2(n764), .I3(n765), .O(n763) );
  INVCKGHD U720 ( .I(n765), .O(n762) );
  INVCKGHD U721 ( .I(n879), .O(n856) );
  ND2HHD U722 ( .I1(n739), .I2(n989), .O(n1001) );
  XNR2HHD U723 ( .I1(n1565), .I2(n821), .O(n989) );
  XNR2KHD U724 ( .I1(n1004), .I2(n1003), .O(n1056) );
  XNR2EHD U725 ( .I1(n1064), .I2(n1063), .O(n1082) );
  INVCHD U726 ( .I(n1062), .O(n1063) );
  ND2HHD U727 ( .I1(n751), .I2(n788), .O(n750) );
  ND3CHD U728 ( .I1(n1050), .I2(n1049), .I3(n1048), .O(n1053) );
  XNR2HHD U729 ( .I1(rnd_25), .I2(n877), .O(n1242) );
  NR2EHD U730 ( .I1(n939), .I2(n938), .O(n940) );
  ND2HHD U731 ( .I1(n701), .I2(n700), .O(n1081) );
  ND2HHD U732 ( .I1(n768), .I2(n1015), .O(n1113) );
  NR2IHD U733 ( .I1(n1061), .I2(n896), .O(n988) );
  NR2EHD U734 ( .I1(rnd_25), .I2(rnd_24), .O(n871) );
  ND3CHD U735 ( .I1(n1306), .I2(n865), .I3(n914), .O(n866) );
  NR2GHD U736 ( .I1(n1167), .I2(n668), .O(n667) );
  ND2DHD U737 ( .I1(n1097), .I2(n1096), .O(n742) );
  ND2DHD U738 ( .I1(n1117), .I2(n1118), .O(n1096) );
  ND2KHD U739 ( .I1(n1306), .I2(n943), .O(n932) );
  ND2DHD U740 ( .I1(n1099), .I2(n1072), .O(n700) );
  INVGHD U741 ( .I(n1140), .O(n991) );
  ND2HHD U742 ( .I1(n889), .I2(n888), .O(n892) );
  ND2HHD U743 ( .I1(n1115), .I2(n1066), .O(n1067) );
  AN3EHD U744 ( .I1(n1305), .I2(n1306), .I3(n1561), .O(n832) );
  NR2GHD U745 ( .I1(rnd_17), .I2(rnd_16), .O(n1305) );
  ND2HHD U746 ( .I1(n1065), .I2(n1252), .O(n1068) );
  XOR2HHD U747 ( .I1(n1207), .I2(n1206), .O(n1205) );
  INVGHD U748 ( .I(n970), .O(n1207) );
  ND3CHD U749 ( .I1(n1561), .I2(n1562), .I3(n1306), .O(n1307) );
  ND2DHD U750 ( .I1(n835), .I2(n1562), .O(n836) );
  ND2DHD U751 ( .I1(n833), .I2(n1562), .O(n837) );
  XOR2HHD U752 ( .I1(n905), .I2(n906), .O(n924) );
  ND2HHD U753 ( .I1(n885), .I2(n886), .O(n905) );
  ND2HHD U754 ( .I1(n1068), .I2(n1067), .O(n1099) );
  INVCHD U755 ( .I(n1105), .O(n1007) );
  ND2DHD U756 ( .I1(n995), .I2(n994), .O(n671) );
  INVCHD U757 ( .I(n1118), .O(n1120) );
  INVCHD U758 ( .I(n1117), .O(n1121) );
  ND2DHD U759 ( .I1(n1214), .I2(n755), .O(n1254) );
  INVKHD U760 ( .I(n1137), .O(n826) );
  INVDHD U761 ( .I(n1144), .O(n1213) );
  XNR2EHD U762 ( .I1(n1252), .I2(n1253), .O(n1263) );
  ND2CHD U763 ( .I1(n1207), .I2(n1206), .O(n1208) );
  INVCHD U764 ( .I(n1233), .O(n1265) );
  ND2CHD U765 ( .I1(n1274), .I2(n1272), .O(n1278) );
  NR2CHD U766 ( .I1(n1274), .I2(n1275), .O(n711) );
  XOR2CHD U767 ( .I1(rkey_next_32), .I2(rkey_next_13), .O(n1453) );
  XOR2CHD U768 ( .I1(rkey_next_1), .I2(rkey_next_36), .O(n1411) );
  XOR2CHD U769 ( .I1(rkey_next_35), .I2(rkey_next_0), .O(n1497) );
  AN3CHD U770 ( .I1(n934), .I2(n1563), .I3(n933), .O(n941) );
  INVCHD U771 ( .I(rnd_23), .O(n767) );
  ND2CHD U772 ( .I1(n937), .I2(n1305), .O(n938) );
  ND2DHD U773 ( .I1(n936), .I2(n935), .O(n939) );
  NR2BHD U774 ( .I1(rnd_5), .I2(rnd_6), .O(n968) );
  XOR2CHD U775 ( .I1(rnd_6), .I2(_keyexpantion_N27 ), .O(n976) );
  ND2DHD U776 ( .I1(n801), .I2(n1568), .O(n1046) );
  AO12EHD U777 ( .B1(n974), .B2(n973), .A1(rnd_16), .O(n993) );
  ND2HHD U778 ( .I1(n977), .I2(_keyexpantion_N27 ), .O(n995) );
  INVCKGHD U779 ( .I(n1242), .O(n882) );
  INVCHD U780 ( .I(n872), .O(n802) );
  ND2CHD U781 ( .I1(n1092), .I2(n1007), .O(n1008) );
  ND2DHD U782 ( .I1(n1005), .I2(n1105), .O(n1006) );
  ND2CHD U783 ( .I1(n1046), .I2(n1044), .O(n1075) );
  XOR2CHD U784 ( .I1(rnd_2), .I2(rnd_7), .O(n972) );
  ND2DHD U785 ( .I1(n1039), .I2(n1038), .O(n1074) );
  XNR2HHD U786 ( .I1(n1558), .I2(n867), .O(n898) );
  NR2EHD U787 ( .I1(n866), .I2(n878), .O(n867) );
  ND2DHD U788 ( .I1(n771), .I2(n977), .O(n952) );
  ND2DHD U789 ( .I1(n952), .I2(n984), .O(n951) );
  NR2CHD U790 ( .I1(n1027), .I2(n753), .O(n798) );
  AN2EHD U791 ( .I1(n753), .I2(n1027), .O(n758) );
  INVDHD U792 ( .I(n1112), .O(n1133) );
  ND2CHD U793 ( .I1(n1113), .I2(n1569), .O(n1116) );
  INVCHD U794 ( .I(n1000), .O(n1002) );
  OA12EHD U795 ( .B1(n983), .B2(n984), .A1(n665), .O(n1004) );
  ND2CHD U796 ( .I1(n1135), .I2(n666), .O(n665) );
  INVCHD U797 ( .I(n1032), .O(n983) );
  XNR3CHD U798 ( .I1(rnd_6), .I2(rnd_16), .I3(n878), .O(n870) );
  XNR2CHD U799 ( .I1(n1203), .I2(n1202), .O(n1245) );
  INVCHD U800 ( .I(n1240), .O(n1203) );
  ND2CHD U801 ( .I1(n1092), .I2(n1091), .O(n1211) );
  AN2CHD U802 ( .I1(n895), .I2(n785), .O(n618) );
  INVCHD U803 ( .I(n1245), .O(n1246) );
  INVCHD U804 ( .I(n1252), .O(n1257) );
  INVCHD U805 ( .I(n1253), .O(n1256) );
  XOR2CHD U806 ( .I1(n1251), .I2(n1250), .O(n1259) );
  OA12EHD U807 ( .B1(n1213), .B2(n1212), .A1(n1211), .O(n1249) );
  INVCHD U808 ( .I(n1210), .O(n1212) );
  OR2CHD U809 ( .I1(n1029), .I2(n1028), .O(n619) );
  ND2CHD U810 ( .I1(n1058), .I2(n1057), .O(n810) );
  INVDHD U811 ( .I(n1273), .O(n712) );
  XNR2CHD U812 ( .I1(n1265), .I2(n1264), .O(n1238) );
  INVCHD U813 ( .I(n1272), .O(n1271) );
  ND2CHD U814 ( .I1(n1579), .I2(rnd_3), .O(n1577) );
  INVCHD U815 ( .I(n943), .O(n1316) );
  NR2BHD U816 ( .I1(rnd_26), .I2(rnd_25), .O(n1311) );
  NR2BHD U817 ( .I1(rnd_12), .I2(rnd_18), .O(n1312) );
  NR2BHD U818 ( .I1(rnd_22), .I2(rnd_29), .O(n1309) );
  NR2BHD U819 ( .I1(rnd_24), .I2(rnd_23), .O(n1310) );
  ND2CHD U820 ( .I1(n1305), .I2(n1568), .O(n1308) );
  INVDHD U821 ( .I(rnd_9), .O(n1555) );
  AN2CHD U822 ( .I1(n1847), .I2(n1846), .O(n1848) );
  ND2CHD U823 ( .I1(n1845), .I2(key_51), .O(n1847) );
  ND2CHD U824 ( .I1(n1807), .I2(Kin_3), .O(n1846) );
  ND2CHD U825 ( .I1(n1852), .I2(rkey_next_3), .O(n1853) );
  MUX2CHD U826 ( .A(n1381), .B(n1380), .S(n1379), .O(n1511) );
  ND2CHD U827 ( .I1(n1845), .I2(key_54), .O(n1831) );
  ND2CHD U828 ( .I1(n1852), .I2(rkey_next_6), .O(n1835) );
  ND2CHD U829 ( .I1(n1851), .I2(key_38), .O(n1836) );
  MUX2CHD U830 ( .A(n1435), .B(n1442), .S(n1434), .O(n1823) );
  ND2CHD U831 ( .I1(n1845), .I2(key_57), .O(n1815) );
  ND2CHD U832 ( .I1(n1852), .I2(rkey_next_9), .O(n1819) );
  ND2CHD U833 ( .I1(n1851), .I2(key_41), .O(n1820) );
  MUX2CHD U834 ( .A(n1424), .B(n1484), .S(n1423), .O(n1806) );
  AN2CHD U835 ( .I1(n1798), .I2(n1797), .O(n1799) );
  ND2CHD U836 ( .I1(n1845), .I2(key_60), .O(n1798) );
  ND2CHD U837 ( .I1(n1807), .I2(Kin_12), .O(n1797) );
  ND2CHD U838 ( .I1(n1852), .I2(rkey_next_12), .O(n1802) );
  MUX2CHD U839 ( .A(n1391), .B(n1390), .S(n1389), .O(n1790) );
  AN2CHD U840 ( .I1(n1782), .I2(n1781), .O(n1783) );
  ND2CHD U841 ( .I1(n1845), .I2(key_63), .O(n1782) );
  ND2CHD U842 ( .I1(n1807), .I2(Kin_15), .O(n1781) );
  ND2CHD U843 ( .I1(n1852), .I2(rkey_next_15), .O(n1786) );
  XNR2CHD U844 ( .I1(n1497), .I2(n1496), .O(n1774) );
  AN2CHD U845 ( .I1(n1766), .I2(n1765), .O(n1767) );
  ND2CHD U846 ( .I1(n1845), .I2(key_50), .O(n1766) );
  ND2CHD U847 ( .I1(n1807), .I2(Kin_2), .O(n1765) );
  ND2CHD U848 ( .I1(n1852), .I2(rkey_next_2), .O(n1770) );
  MUX2CHD U849 ( .A(n1352), .B(n1412), .S(n1351), .O(n1758) );
  ND2CHD U850 ( .I1(n1845), .I2(key_53), .O(n1750) );
  ND2CHD U851 ( .I1(n1852), .I2(rkey_next_5), .O(n1754) );
  ND2CHD U852 ( .I1(n1851), .I2(key_37), .O(n1755) );
  MUX2CHD U853 ( .A(n1444), .B(n1462), .S(n1443), .O(n1742) );
  AN2CHD U854 ( .I1(n1734), .I2(n1733), .O(n1735) );
  ND2CHD U855 ( .I1(n1845), .I2(key_56), .O(n1734) );
  ND2CHD U856 ( .I1(n1807), .I2(Kin_8), .O(n1733) );
  ND2CHD U857 ( .I1(n1852), .I2(rkey_next_8), .O(n1738) );
  MUX2CHD U858 ( .A(n1487), .B(n1486), .S(n1485), .O(n1726) );
  ND2CHD U859 ( .I1(n1845), .I2(key_59), .O(n1718) );
  ND2CHD U860 ( .I1(n1852), .I2(rkey_next_11), .O(n1722) );
  ND2CHD U861 ( .I1(n1851), .I2(key_43), .O(n1723) );
  MUX2CHD U862 ( .A(n1361), .B(n1400), .S(n1360), .O(n1710) );
  ND2CHD U863 ( .I1(n1845), .I2(key_62), .O(n1702) );
  ND2CHD U864 ( .I1(n1852), .I2(rkey_next_14), .O(n1706) );
  ND2CHD U865 ( .I1(n1851), .I2(key_46), .O(n1707) );
  MUX2CHD U866 ( .A(n1475), .B(n1474), .S(n1473), .O(n1694) );
  ND2CHD U867 ( .I1(n1845), .I2(key_49), .O(n1686) );
  ND2CHD U868 ( .I1(n1852), .I2(rkey_next_1), .O(n1690) );
  ND2CHD U869 ( .I1(n1851), .I2(key_33), .O(n1691) );
  XNR2CHD U870 ( .I1(n1414), .I2(n1413), .O(n1682) );
  MUX2CHD U871 ( .A(rkey_1), .B(n1689), .S(n1412), .O(n1413) );
  ND2CHD U872 ( .I1(n1845), .I2(key_52), .O(n1674) );
  ND2CHD U873 ( .I1(n1852), .I2(rkey_next_4), .O(n1678) );
  ND2CHD U874 ( .I1(n1851), .I2(key_36), .O(n1679) );
  MUX2CHD U875 ( .A(n1465), .B(n1464), .S(n1463), .O(n1506) );
  AN2CHD U876 ( .I1(n1661), .I2(n1660), .O(n1662) );
  ND2CHD U877 ( .I1(n1845), .I2(key_55), .O(n1661) );
  ND2CHD U878 ( .I1(n1807), .I2(Kin_7), .O(n1660) );
  ND2CHD U879 ( .I1(n1852), .I2(rkey_next_7), .O(n1665) );
  MUX2CHD U880 ( .A(n1371), .B(n1433), .S(n1370), .O(n1653) );
  ND2CHD U881 ( .I1(n1845), .I2(key_58), .O(n1645) );
  ND2CHD U882 ( .I1(n1852), .I2(rkey_next_10), .O(n1649) );
  ND2CHD U883 ( .I1(n1851), .I2(key_42), .O(n1650) );
  MUX2CHD U884 ( .A(n1402), .B(n1422), .S(n1401), .O(n1637) );
  AN2CHD U885 ( .I1(n1629), .I2(n1628), .O(n1630) );
  ND2CHD U886 ( .I1(n1845), .I2(key_61), .O(n1629) );
  ND2CHD U887 ( .I1(n1807), .I2(Kin_13), .O(n1628) );
  ND2CHD U888 ( .I1(n1852), .I2(rkey_next_13), .O(n1633) );
  ND2CHD U889 ( .I1(n1807), .I2(Kin_29), .O(n1624) );
  XNR2CHD U890 ( .I1(n1453), .I2(n1452), .O(n1621) );
  MUX2CHD U891 ( .A(rkey_13), .B(n1632), .S(n1474), .O(n1452) );
  XNR3CHD U892 ( .I1(rkey_0), .I2(n1411), .I3(n1497), .O(n1548) );
  ND2CHD U893 ( .I1(n1807), .I2(Kin_48), .O(n1587) );
  INVCHD U894 ( .I(n1852), .O(n1551) );
  INVCHD U895 ( .I(n915), .O(n854) );
  ND2CHD U896 ( .I1(n844), .I2(n843), .O(n846) );
  INVCHD U897 ( .I(rnd_4), .O(n843) );
  INVDHD U898 ( .I(n990), .O(n740) );
  ND2DHD U899 ( .I1(n990), .I2(n788), .O(n739) );
  NR2EHD U900 ( .I1(n869), .I2(n868), .O(n973) );
  INVCHD U901 ( .I(n1039), .O(n887) );
  INVDHD U902 ( .I(n1251), .O(n889) );
  ND2CHD U903 ( .I1(n969), .I2(n1579), .O(n1037) );
  ND2CHD U904 ( .I1(n1013), .I2(n863), .O(n874) );
  NR2BHD U905 ( .I1(n828), .I2(n830), .O(n829) );
  ND2CHD U906 ( .I1(n943), .I2(rnd_20), .O(n828) );
  INVCHD U907 ( .I(n830), .O(n831) );
  NR2BHD U908 ( .I1(rnd_8), .I2(rnd_7), .O(n853) );
  AN2CHD U909 ( .I1(n941), .I2(n767), .O(n625) );
  ND2CHD U910 ( .I1(n745), .I2(n1579), .O(n1105) );
  INVCHD U911 ( .I(n985), .O(n986) );
  INVCHD U912 ( .I(n1044), .O(n1090) );
  XNR2CHD U913 ( .I1(n1579), .I2(n981), .O(n1108) );
  XOR2CHD U914 ( .I1(rnd_13), .I2(rnd_3), .O(n981) );
  ND2DHD U915 ( .I1(n823), .I2(n790), .O(n789) );
  AN2CHD U916 ( .I1(n934), .I2(n1562), .O(n790) );
  INVCHD U917 ( .I(n822), .O(n823) );
  ND2DHD U918 ( .I1(n786), .I2(n974), .O(n751) );
  AN2CHD U919 ( .I1(n974), .I2(n824), .O(n749) );
  INVCHD U920 ( .I(n1073), .O(n1098) );
  ND2CHD U921 ( .I1(n1071), .I2(n1070), .O(n1100) );
  ND2CHD U922 ( .I1(n1069), .I2(rnd_14), .O(n1070) );
  INVCHD U923 ( .I(n993), .O(n992) );
  AN2CHD U924 ( .I1(n1106), .I2(n1105), .O(n1112) );
  ND2DHD U925 ( .I1(n1136), .I2(rnd_12), .O(n1106) );
  AN2CHD U926 ( .I1(n1001), .I2(n998), .O(n622) );
  ND2DHD U927 ( .I1(n1052), .I2(n1054), .O(n697) );
  INVCHD U928 ( .I(n1076), .O(n1049) );
  ND2CHD U929 ( .I1(n1077), .I2(n1075), .O(n1050) );
  ND2DHD U930 ( .I1(n673), .I2(n669), .O(n698) );
  ND2CHD U931 ( .I1(n884), .I2(rnd_30), .O(n885) );
  ND2CHD U932 ( .I1(n1039), .I2(n1045), .O(n891) );
  ND2CHD U933 ( .I1(n887), .I2(n1090), .O(n888) );
  ND2DHD U934 ( .I1(n1140), .I2(n912), .O(n911) );
  XNR2CHD U935 ( .I1(rnd_5), .I2(n1037), .O(n1038) );
  NR2BHD U936 ( .I1(rnd_14), .I2(n869), .O(n839) );
  ND2CHD U937 ( .I1(n853), .I2(n914), .O(n879) );
  INVCHD U938 ( .I(n910), .O(n851) );
  XNR2HHD U939 ( .I1(rnd_8), .I2(n944), .O(n982) );
  NR2CHD U940 ( .I1(n1014), .I2(n1033), .O(n1015) );
  XOR2EHD U941 ( .I1(rnd_28), .I2(n949), .O(n970) );
  ND2DHD U942 ( .I1(n768), .I2(n948), .O(n949) );
  NR2CHD U943 ( .I1(n947), .I2(n1033), .O(n948) );
  XNR2CHD U944 ( .I1(rnd_7), .I2(n971), .O(n950) );
  ND2DHD U945 ( .I1(n691), .I2(n1023), .O(n690) );
  XNR2CHD U946 ( .I1(rnd_31), .I2(n1061), .O(n1064) );
  ND2DHD U947 ( .I1(n702), .I2(n1100), .O(n701) );
  ND3CHD U948 ( .I1(n1068), .I2(n1067), .I3(n703), .O(n702) );
  INVCKGHD U949 ( .I(n1111), .O(n1131) );
  OR2CHD U950 ( .I1(n754), .I2(n982), .O(n621) );
  INVCHD U951 ( .I(n1107), .O(n754) );
  NR2CHD U952 ( .I1(n788), .I2(n789), .O(n787) );
  ND2DHD U953 ( .I1(n1073), .I2(rnd_25), .O(n719) );
  INVDHD U954 ( .I(n1078), .O(n645) );
  INVDHD U955 ( .I(n1024), .O(n893) );
  ND2CHD U956 ( .I1(n903), .I2(n902), .O(n904) );
  INVCHD U957 ( .I(n906), .O(n903) );
  INVCHD U958 ( .I(n905), .O(n902) );
  XNR3CHD U959 ( .I1(n1061), .I2(n897), .I3(n896), .O(n923) );
  ND2CHD U960 ( .I1(n906), .I2(n905), .O(n925) );
  ND2DHD U961 ( .I1(n913), .I2(n991), .O(n638) );
  ND2DHD U962 ( .I1(n911), .I2(n989), .O(n637) );
  INVCHD U963 ( .I(n912), .O(n913) );
  ND3CHD U964 ( .I1(n974), .I2(n824), .I3(n1350), .O(n678) );
  XNR2CHD U965 ( .I1(n982), .I2(n1214), .O(n1210) );
  MAO222CHD U966 ( .A1(n1135), .B1(n950), .C1(rnd_17), .O(n1206) );
  ND2CHD U967 ( .I1(n1110), .I2(n953), .O(n954) );
  INVCHD U968 ( .I(n952), .O(n953) );
  XOR2EHD U969 ( .I1(n1205), .I2(n1204), .O(n1199) );
  INVDHD U970 ( .I(n1159), .O(n687) );
  ND2DHD U971 ( .I1(n1165), .I2(n733), .O(n686) );
  ND2CHD U972 ( .I1(n1163), .I2(n1162), .O(n1165) );
  INVCHD U973 ( .I(n1161), .O(n1162) );
  XNR2EHD U974 ( .I1(n923), .I2(n924), .O(n1167) );
  ND2DHD U975 ( .I1(n1166), .I2(_keyexpantion_N27 ), .O(n1171) );
  ND2DHD U976 ( .I1(n806), .I2(n805), .O(n1166) );
  ND2CHD U977 ( .I1(n1102), .I2(n1101), .O(n1103) );
  ND2CHD U978 ( .I1(n1127), .I2(n1128), .O(n1104) );
  XOR2CHD U979 ( .I1(n1134), .I2(n616), .O(n1147) );
  MAO222CHD U980 ( .A1(n1131), .B1(n1130), .C1(n1110), .O(n1134) );
  XOR2CHD U981 ( .I1(n1133), .I2(n1132), .O(n616) );
  XOR2CHD U982 ( .I1(n1213), .I2(rnd_28), .O(n1145) );
  MAO222CHD U983 ( .A1(n1143), .B1(n1142), .C1(n1141), .O(n1146) );
  XNR2CHD U984 ( .I1(n1136), .I2(n1135), .O(n1142) );
  MAO222CHD U985 ( .A1(n1140), .B1(n1139), .C1(n1138), .O(n1141) );
  ND2CHD U986 ( .I1(n1137), .I2(_keyexpantion_N26 ), .O(n1139) );
  OA12EHD U987 ( .B1(n1126), .B2(n1129), .A1(n1125), .O(n1149) );
  INVCHD U988 ( .I(n1122), .O(n1124) );
  OR2CHD U989 ( .I1(n1004), .I2(n1003), .O(n815) );
  ND2CHD U990 ( .I1(n900), .I2(n899), .O(n901) );
  INVCHD U991 ( .I(n956), .O(n929) );
  ND2DHD U992 ( .I1(n926), .I2(n925), .O(n962) );
  ND2CHD U993 ( .I1(n924), .I2(n923), .O(n926) );
  OA12EHD U994 ( .B1(n929), .B2(n961), .A1(n960), .O(n1195) );
  ND2CHD U995 ( .I1(n959), .I2(n958), .O(n960) );
  INVCHD U996 ( .I(n957), .O(n958) );
  XNR2CHD U997 ( .I1(rnd_3), .I2(rnd_2), .O(n1190) );
  INVCHD U998 ( .I(n716), .O(n715) );
  XNR3CHD U999 ( .I1(n1262), .I2(n1261), .I3(n1260), .O(n1267) );
  XOR2CHD U1000 ( .I1(n1244), .I2(n1243), .O(n1262) );
  XNR2CHD U1001 ( .I1(n1234), .I2(n1233), .O(n1217) );
  INVCHD U1002 ( .I(n1235), .O(n1237) );
  ND2HHD U1003 ( .I1(n775), .I2(n774), .O(n1177) );
  INVDHD U1004 ( .I(n1169), .O(n774) );
  INVDHD U1005 ( .I(n1168), .O(n775) );
  INVCHD U1006 ( .I(n1183), .O(n1175) );
  INVDHD U1007 ( .I(n964), .O(n967) );
  NR2BHD U1008 ( .I1(n657), .I2(n1059), .O(n811) );
  ND2HHD U1009 ( .I1(n965), .I2(n964), .O(n1230) );
  INVCHD U1010 ( .I(n1285), .O(n1280) );
  INVCHD U1011 ( .I(sel), .O(n1294) );
  ND3CHD U1012 ( .I1(n712), .I2(n1277), .I3(n711), .O(n710) );
  INVCHD U1013 ( .I(Krdy), .O(n1327) );
  XOR2CHD U1014 ( .I1(n818), .I2(n1548), .O(n626) );
  OR2CHD U1015 ( .I1(Drdy), .I2(n1297), .O(n1298) );
  INVCHD U1016 ( .I(rnd_30), .O(n1568) );
  INVCHD U1017 ( .I(rnd_29), .O(n1569) );
  INVCHD U1018 ( .I(rnd_26), .O(n1565) );
  INVDHD U1019 ( .I(rnd_25), .O(n1566) );
  INVDHD U1020 ( .I(rnd_24), .O(n1564) );
  INVDHD U1021 ( .I(rnd_22), .O(n1563) );
  INVCHD U1022 ( .I(rnd_21), .O(n788) );
  INVDHD U1023 ( .I(rnd_18), .O(n1560) );
  INVDHD U1024 ( .I(rnd_16), .O(n909) );
  INVCHD U1025 ( .I(rnd_12), .O(n1557) );
  INVDHD U1026 ( .I(rnd_11), .O(n1558) );
  INVDHD U1027 ( .I(rnd_10), .O(n1556) );
  INVCHD U1028 ( .I(Drdy), .O(n1348) );
  ND2CHD U1029 ( .I1(n1807), .I2(Kin_35), .O(n1613) );
  ND2CHD U1030 ( .I1(n1807), .I2(Kin_38), .O(n1607) );
  ND2CHD U1031 ( .I1(n1807), .I2(Kin_41), .O(n1601) );
  ND2CHD U1032 ( .I1(n1807), .I2(Kin_44), .O(n1595) );
  ND2CHD U1033 ( .I1(n1807), .I2(Kin_47), .O(n1589) );
  ND2CHD U1034 ( .I1(n1807), .I2(Kin_34), .O(n1615) );
  ND2CHD U1035 ( .I1(n1807), .I2(Kin_37), .O(n1609) );
  ND2CHD U1036 ( .I1(n1807), .I2(Kin_40), .O(n1603) );
  ND2CHD U1037 ( .I1(n1807), .I2(Kin_43), .O(n1597) );
  ND2CHD U1038 ( .I1(n1807), .I2(Kin_46), .O(n1591) );
  ND2CHD U1039 ( .I1(n1807), .I2(Kin_33), .O(n1617) );
  ND2CHD U1040 ( .I1(n1807), .I2(Kin_36), .O(n1611) );
  ND2CHD U1041 ( .I1(n1807), .I2(Kin_39), .O(n1605) );
  ND2CHD U1042 ( .I1(n1807), .I2(Kin_42), .O(n1599) );
  ND2CHD U1043 ( .I1(n1807), .I2(Kin_45), .O(n1593) );
  NR2BHD U1044 ( .I1(n1578), .I2(n1329), .O(n1330) );
  ND2CHD U1045 ( .I1(n1807), .I2(Kin_32), .O(n1619) );
  NR2BHD U1046 ( .I1(Drdy), .I2(rnd_13), .O(n1301) );
  NR2BHD U1047 ( .I1(rnd_21), .I2(rnd_27), .O(n1304) );
  NR2BHD U1048 ( .I1(n1316), .I2(n1315), .O(n1317) );
  ND2CHD U1049 ( .I1(n1326), .I2(n1325), .O(n611) );
  AO222CHD U1050 ( .A1(n1571), .A2(Dout_6), .B1(n1573), .B2(Din_6), .C1(n1572), .C2(dat_next_6), .O(n510) );
  ND2CHD U1051 ( .I1(n1441), .I2(n1440), .O(n494) );
  AO222CHD U1052 ( .A1(n1571), .A2(Dout_5), .B1(n1573), .B2(Din_5), .C1(n1572), .C2(dat_next_5), .O(n511) );
  ND2CHD U1053 ( .I1(n1451), .I2(n1450), .O(n495) );
  AO222CHD U1054 ( .A1(n1571), .A2(Dout_13), .B1(n1573), .B2(Din_13), .C1(n1572), .C2(dat_next_13), .O(n503) );
  ND2CHD U1055 ( .I1(n1461), .I2(n1460), .O(n487) );
  AO222CHD U1056 ( .A1(n1571), .A2(Dout_4), .B1(n1573), .B2(Din_4), .C1(n1572), .C2(dat_next_4), .O(n512) );
  ND2CHD U1057 ( .I1(n1472), .I2(n1471), .O(n496) );
  AO222CHD U1058 ( .A1(n1571), .A2(Dout_3), .B1(n1573), .B2(Din_3), .C1(n1572), .C2(dat_next_3), .O(n513) );
  ND2CHD U1059 ( .I1(n1388), .I2(n1387), .O(n497) );
  AO222CHD U1060 ( .A1(n1571), .A2(Dout_11), .B1(n1573), .B2(Din_11), .C1(n1572), .C2(dat_next_11), .O(n505) );
  ND2CHD U1061 ( .I1(n1369), .I2(n1368), .O(n489) );
  AO222CHD U1062 ( .A1(n1571), .A2(Dout_2), .B1(n1573), .B2(Din_2), .C1(n1572), .C2(dat_next_2), .O(n514) );
  ND2CHD U1063 ( .I1(n1359), .I2(n1358), .O(n498) );
  AO222CHD U1064 ( .A1(n1571), .A2(Dout_1), .B1(n1573), .B2(Din_1), .C1(n1572), .C2(dat_next_1), .O(n515) );
  ND2CHD U1065 ( .I1(n1421), .I2(n1420), .O(n499) );
  AO222CHD U1066 ( .A1(n1571), .A2(Dout_9), .B1(n1573), .B2(Din_9), .C1(n1572), .C2(dat_next_9), .O(n507) );
  ND2CHD U1067 ( .I1(n1432), .I2(n1431), .O(n491) );
  AO222CHD U1068 ( .A1(n1571), .A2(Dout_7), .B1(n1573), .B2(Din_7), .C1(n1572), .C2(dat_next_7), .O(n509) );
  ND2CHD U1069 ( .I1(n1378), .I2(n1377), .O(n493) );
  AO222CHD U1070 ( .A1(n1571), .A2(Dout_15), .B1(n1573), .B2(Din_15), .C1(n1572), .C2(dat_next_15), .O(n501) );
  ND2CHD U1071 ( .I1(n1505), .I2(n1504), .O(n484) );
  AO222CHD U1072 ( .A1(n1571), .A2(Dout_14), .B1(n1573), .B2(Din_14), .C1(n1572), .C2(dat_next_14), .O(n502) );
  ND2CHD U1073 ( .I1(n1483), .I2(n1482), .O(n486) );
  AO222CHD U1074 ( .A1(n1571), .A2(Dout_12), .B1(n1573), .B2(Din_12), .C1(n1572), .C2(dat_next_12), .O(n504) );
  ND2CHD U1075 ( .I1(n1399), .I2(n1398), .O(n488) );
  AO222CHD U1076 ( .A1(n1571), .A2(Dout_10), .B1(n1573), .B2(Din_10), .C1(n1572), .C2(dat_next_10), .O(n506) );
  ND2CHD U1077 ( .I1(n1410), .I2(n1409), .O(n490) );
  AO222CHD U1078 ( .A1(n1571), .A2(Dout_8), .B1(n1573), .B2(Din_8), .C1(n1572), .C2(dat_next_8), .O(n508) );
  ND2CHD U1079 ( .I1(n1494), .I2(n1493), .O(n492) );
  ND2CHD U1080 ( .I1(n1572), .I2(dat_next_0), .O(n1575) );
  ND2CHD U1081 ( .I1(n1571), .I2(Dout_0), .O(n1576) );
  MUX2CHD U1082 ( .A(key_0), .B(Kin_0), .S(n1807), .O(n517) );
  MUX2CHD U1083 ( .A(key_1), .B(Kin_1), .S(n1807), .O(n518) );
  MUX2CHD U1084 ( .A(key_2), .B(Kin_2), .S(n1807), .O(n519) );
  MUX2CHD U1085 ( .A(key_3), .B(Kin_3), .S(n1807), .O(n520) );
  MUX2CHD U1086 ( .A(key_4), .B(Kin_4), .S(n1807), .O(n521) );
  MUX2CHD U1087 ( .A(key_5), .B(Kin_5), .S(n1807), .O(n522) );
  MUX2CHD U1088 ( .A(key_6), .B(Kin_6), .S(n1807), .O(n523) );
  MUX2CHD U1089 ( .A(key_7), .B(Kin_7), .S(n1807), .O(n524) );
  MUX2CHD U1090 ( .A(key_8), .B(Kin_8), .S(n1807), .O(n525) );
  MUX2CHD U1091 ( .A(key_9), .B(Kin_9), .S(n1807), .O(n526) );
  MUX2CHD U1092 ( .A(key_10), .B(Kin_10), .S(n1807), .O(n527) );
  MUX2CHD U1093 ( .A(key_11), .B(Kin_11), .S(n1807), .O(n528) );
  MUX2CHD U1094 ( .A(key_12), .B(Kin_12), .S(n1807), .O(n529) );
  MUX2CHD U1095 ( .A(key_13), .B(Kin_13), .S(n1807), .O(n530) );
  MUX2CHD U1096 ( .A(key_14), .B(Kin_14), .S(n1807), .O(n531) );
  MUX2CHD U1097 ( .A(key_15), .B(Kin_15), .S(n1807), .O(n532) );
  MUX2CHD U1098 ( .A(key_16), .B(Kin_16), .S(n1807), .O(n533) );
  MUX2CHD U1099 ( .A(key_17), .B(Kin_17), .S(n1807), .O(n534) );
  MUX2CHD U1100 ( .A(key_18), .B(Kin_18), .S(n1807), .O(n535) );
  MUX2CHD U1101 ( .A(key_19), .B(Kin_19), .S(n1807), .O(n536) );
  MUX2CHD U1102 ( .A(key_20), .B(Kin_20), .S(n1807), .O(n537) );
  MUX2CHD U1103 ( .A(key_21), .B(Kin_21), .S(n1807), .O(n538) );
  MUX2CHD U1104 ( .A(key_22), .B(Kin_22), .S(n1807), .O(n539) );
  MUX2CHD U1105 ( .A(key_23), .B(Kin_23), .S(n1807), .O(n540) );
  MUX2CHD U1106 ( .A(key_24), .B(Kin_24), .S(n1807), .O(n541) );
  MUX2CHD U1107 ( .A(key_25), .B(Kin_25), .S(n1807), .O(n542) );
  MUX2CHD U1108 ( .A(key_26), .B(Kin_26), .S(n1807), .O(n543) );
  MUX2CHD U1109 ( .A(key_27), .B(Kin_27), .S(n1807), .O(n544) );
  MUX2CHD U1110 ( .A(key_28), .B(Kin_28), .S(n1807), .O(n545) );
  MUX2CHD U1111 ( .A(key_29), .B(Kin_29), .S(n1807), .O(n546) );
  MUX2CHD U1112 ( .A(key_30), .B(Kin_30), .S(n1807), .O(n547) );
  MUX2CHD U1113 ( .A(key_31), .B(Kin_31), .S(n1807), .O(n548) );
  MUX2CHD U1114 ( .A(key_49), .B(Kin_49), .S(n1807), .O(n566) );
  MUX2CHD U1115 ( .A(key_50), .B(Kin_50), .S(n1807), .O(n567) );
  MUX2CHD U1116 ( .A(key_51), .B(Kin_51), .S(n1807), .O(n568) );
  MUX2CHD U1117 ( .A(key_52), .B(Kin_52), .S(n1807), .O(n569) );
  MUX2CHD U1118 ( .A(key_53), .B(Kin_53), .S(n1807), .O(n570) );
  MUX2CHD U1119 ( .A(key_54), .B(Kin_54), .S(n1807), .O(n571) );
  MUX2CHD U1120 ( .A(key_55), .B(Kin_55), .S(n1807), .O(n572) );
  MUX2CHD U1121 ( .A(key_56), .B(Kin_56), .S(n1807), .O(n573) );
  MUX2CHD U1122 ( .A(key_57), .B(Kin_57), .S(n1807), .O(n574) );
  MUX2CHD U1123 ( .A(key_58), .B(Kin_58), .S(n1807), .O(n575) );
  MUX2CHD U1124 ( .A(key_59), .B(Kin_59), .S(n1807), .O(n576) );
  MUX2CHD U1125 ( .A(key_60), .B(Kin_60), .S(n1807), .O(n577) );
  MUX2CHD U1126 ( .A(key_61), .B(Kin_61), .S(n1807), .O(n578) );
  MUX2CHD U1127 ( .A(key_62), .B(Kin_62), .S(n1807), .O(n579) );
  MUX2CHD U1128 ( .A(key_63), .B(Kin_63), .S(n1807), .O(n580) );
  MUX2CHD U1129 ( .A(rnd_30), .B(rnd_31), .S(n1570), .O(n612) );
  MUX2CHD U1130 ( .A(rnd_27), .B(rnd_28), .S(n1570), .O(n583) );
  MUX2CHD U1131 ( .A(rnd_26), .B(rnd_27), .S(n1570), .O(n584) );
  MUX2CHD U1132 ( .A(rnd_23), .B(rnd_24), .S(n1570), .O(n587) );
  MUX2CHD U1133 ( .A(rnd_22), .B(rnd_23), .S(n1570), .O(n588) );
  MXL2CHD U1134 ( .A(n1562), .B(n788), .S(n1570), .OB(n590) );
  MUX2CHD U1135 ( .A(rnd_17), .B(rnd_18), .S(n1570), .O(n593) );
  MUX2CHD U1136 ( .A(rnd_16), .B(rnd_17), .S(n1570), .O(n594) );
  MUX2CHD U1137 ( .A(rnd_13), .B(rnd_14), .S(n1570), .O(n597) );
  MUX2CHD U1138 ( .A(rnd_12), .B(rnd_13), .S(n1570), .O(n598) );
  INVCHD U1139 ( .I(rnd_8), .O(n1554) );
  MUX2CHD U1140 ( .A(rnd_7), .B(rnd_8), .S(n1570), .O(n603) );
  MUX2CHD U1141 ( .A(rnd_6), .B(rnd_7), .S(n1570), .O(n604) );
  MUX2CHD U1142 ( .A(rnd_5), .B(rnd_6), .S(n1570), .O(n605) );
  MUX2CHD U1143 ( .A(rnd_4), .B(rnd_5), .S(n1570), .O(n606) );
  MUX2CHD U1144 ( .A(rnd_3), .B(rnd_4), .S(n1570), .O(n607) );
  MUX2CHD U1145 ( .A(rnd_2), .B(rnd_3), .S(n1570), .O(n608) );
  AN2CHD U1146 ( .I1(n1854), .I2(n1853), .O(n1855) );
  ND2CHD U1147 ( .I1(n1851), .I2(key_35), .O(n1854) );
  AN2CHD U1148 ( .I1(n1840), .I2(n1839), .O(n1841) );
  ND2CHD U1149 ( .I1(n1852), .I2(rkey_next_19), .O(n1840) );
  ND2CHD U1150 ( .I1(n1807), .I2(Kin_19), .O(n1839) );
  ND2CHD U1151 ( .I1(n1335), .I2(n1613), .O(n418) );
  AN2CHD U1152 ( .I1(n1334), .I2(n1333), .O(n1335) );
  ND2CHD U1153 ( .I1(rkey_next_19), .I2(n1584), .O(n1333) );
  ND2CHD U1154 ( .I1(n1852), .I2(rkey_next_35), .O(n1334) );
  ND2CHD U1155 ( .I1(n1513), .I2(n1512), .O(n419) );
  ND2CHD U1156 ( .I1(n1511), .I2(n1852), .O(n1513) );
  AN2CHD U1157 ( .I1(n1836), .I2(n1835), .O(n1837) );
  AN2CHD U1158 ( .I1(n1831), .I2(n1830), .O(n1832) );
  AN2CHD U1159 ( .I1(n1827), .I2(n1826), .O(n1828) );
  ND2CHD U1160 ( .I1(n1807), .I2(Kin_22), .O(n1826) );
  ND2CHD U1161 ( .I1(n1852), .I2(rkey_next_22), .O(n1827) );
  ND2CHD U1162 ( .I1(n1528), .I2(n1607), .O(n422) );
  AN2CHD U1163 ( .I1(n1527), .I2(n1526), .O(n1528) );
  ND2CHD U1164 ( .I1(rkey_next_22), .I2(n1584), .O(n1526) );
  ND2CHD U1165 ( .I1(n1852), .I2(rkey_next_38), .O(n1527) );
  AN2CHD U1166 ( .I1(n1820), .I2(n1819), .O(n1821) );
  AN2CHD U1167 ( .I1(n1815), .I2(n1814), .O(n1816) );
  AN2CHD U1168 ( .I1(n1811), .I2(n1810), .O(n1812) );
  ND2CHD U1169 ( .I1(n1852), .I2(rkey_next_25), .O(n1811) );
  ND2CHD U1170 ( .I1(n1807), .I2(Kin_25), .O(n1810) );
  ND2CHD U1171 ( .I1(n1534), .I2(n1601), .O(n426) );
  AN2CHD U1172 ( .I1(n1533), .I2(n1532), .O(n1534) );
  ND2CHD U1173 ( .I1(rkey_next_25), .I2(n1584), .O(n1532) );
  ND2CHD U1174 ( .I1(n1852), .I2(rkey_next_41), .O(n1533) );
  AN2CHD U1175 ( .I1(n1803), .I2(n1802), .O(n1804) );
  ND2CHD U1176 ( .I1(n1851), .I2(key_44), .O(n1803) );
  AN2CHD U1177 ( .I1(n1794), .I2(n1793), .O(n1795) );
  ND2CHD U1178 ( .I1(n1807), .I2(Kin_28), .O(n1793) );
  ND2CHD U1179 ( .I1(n1852), .I2(rkey_next_28), .O(n1794) );
  ND2CHD U1180 ( .I1(n1341), .I2(n1595), .O(n430) );
  AN2CHD U1181 ( .I1(n1340), .I2(n1339), .O(n1341) );
  ND2CHD U1182 ( .I1(rkey_next_28), .I2(n1584), .O(n1339) );
  ND2CHD U1183 ( .I1(n1852), .I2(rkey_next_44), .O(n1340) );
  AN2CHD U1184 ( .I1(n1787), .I2(n1786), .O(n1788) );
  ND2CHD U1185 ( .I1(n1851), .I2(key_47), .O(n1787) );
  AN2CHD U1186 ( .I1(n1778), .I2(n1777), .O(n1779) );
  ND2CHD U1187 ( .I1(n1807), .I2(Kin_31), .O(n1777) );
  ND2CHD U1188 ( .I1(n1852), .I2(rkey_next_31), .O(n1778) );
  ND2CHD U1189 ( .I1(n1531), .I2(n1589), .O(n434) );
  AN2CHD U1190 ( .I1(n1530), .I2(n1529), .O(n1531) );
  ND2CHD U1191 ( .I1(rkey_next_31), .I2(n1584), .O(n1529) );
  ND2CHD U1192 ( .I1(n1852), .I2(rkey_next_47), .O(n1530) );
  AN2CHD U1193 ( .I1(n1771), .I2(n1770), .O(n1772) );
  ND2CHD U1194 ( .I1(n1851), .I2(key_34), .O(n1771) );
  AN2CHD U1195 ( .I1(n1762), .I2(n1761), .O(n1763) );
  ND2CHD U1196 ( .I1(n1807), .I2(Kin_18), .O(n1761) );
  ND2CHD U1197 ( .I1(n1852), .I2(rkey_next_18), .O(n1762) );
  ND2CHD U1198 ( .I1(n1338), .I2(n1615), .O(n438) );
  AN2CHD U1199 ( .I1(n1337), .I2(n1336), .O(n1338) );
  ND2CHD U1200 ( .I1(rkey_next_18), .I2(n1584), .O(n1336) );
  ND2CHD U1201 ( .I1(n1852), .I2(rkey_next_34), .O(n1337) );
  AN2CHD U1202 ( .I1(n1755), .I2(n1754), .O(n1756) );
  AN2CHD U1203 ( .I1(n1750), .I2(n1749), .O(n1751) );
  AN2CHD U1204 ( .I1(n1746), .I2(n1745), .O(n1747) );
  ND2CHD U1205 ( .I1(n1807), .I2(Kin_21), .O(n1745) );
  ND2CHD U1206 ( .I1(n1852), .I2(rkey_next_21), .O(n1746) );
  ND2CHD U1207 ( .I1(n1522), .I2(n1609), .O(n442) );
  AN2CHD U1208 ( .I1(n1521), .I2(n1520), .O(n1522) );
  ND2CHD U1209 ( .I1(rkey_next_21), .I2(n1584), .O(n1520) );
  ND2CHD U1210 ( .I1(n1852), .I2(rkey_next_37), .O(n1521) );
  AN2CHD U1211 ( .I1(n1739), .I2(n1738), .O(n1740) );
  ND2CHD U1212 ( .I1(n1851), .I2(key_40), .O(n1739) );
  AN2CHD U1213 ( .I1(n1730), .I2(n1729), .O(n1731) );
  ND2CHD U1214 ( .I1(n1852), .I2(rkey_next_24), .O(n1730) );
  ND2CHD U1215 ( .I1(n1807), .I2(Kin_24), .O(n1729) );
  ND2CHD U1216 ( .I1(n1537), .I2(n1603), .O(n446) );
  AN2CHD U1217 ( .I1(n1536), .I2(n1535), .O(n1537) );
  ND2CHD U1218 ( .I1(rkey_next_24), .I2(n1584), .O(n1535) );
  ND2CHD U1219 ( .I1(n1852), .I2(rkey_next_40), .O(n1536) );
  AN2CHD U1220 ( .I1(n1723), .I2(n1722), .O(n1724) );
  AN2CHD U1221 ( .I1(n1718), .I2(n1717), .O(n1719) );
  AN2CHD U1222 ( .I1(n1714), .I2(n1713), .O(n1715) );
  ND2CHD U1223 ( .I1(n1807), .I2(Kin_27), .O(n1713) );
  ND2CHD U1224 ( .I1(n1852), .I2(rkey_next_27), .O(n1714) );
  ND2CHD U1225 ( .I1(n1344), .I2(n1597), .O(n450) );
  AN2CHD U1226 ( .I1(n1343), .I2(n1342), .O(n1344) );
  ND2CHD U1227 ( .I1(rkey_next_27), .I2(n1584), .O(n1342) );
  ND2CHD U1228 ( .I1(n1852), .I2(rkey_next_43), .O(n1343) );
  AN2CHD U1229 ( .I1(n1707), .I2(n1706), .O(n1708) );
  AN2CHD U1230 ( .I1(n1702), .I2(n1701), .O(n1703) );
  AN2CHD U1231 ( .I1(n1698), .I2(n1697), .O(n1699) );
  ND2CHD U1232 ( .I1(n1852), .I2(rkey_next_30), .O(n1698) );
  ND2CHD U1233 ( .I1(n1807), .I2(Kin_30), .O(n1697) );
  ND2CHD U1234 ( .I1(n1519), .I2(n1591), .O(n454) );
  AN2CHD U1235 ( .I1(n1518), .I2(n1517), .O(n1519) );
  ND2CHD U1236 ( .I1(rkey_next_30), .I2(n1584), .O(n1517) );
  ND2CHD U1237 ( .I1(n1852), .I2(rkey_next_46), .O(n1518) );
  AN2CHD U1238 ( .I1(n1691), .I2(n1690), .O(n1692) );
  AN2CHD U1239 ( .I1(n1686), .I2(n1685), .O(n1687) );
  ND2CHD U1240 ( .I1(n1332), .I2(n1331), .O(n457) );
  ND2CHD U1241 ( .I1(n1852), .I2(rkey_next_17), .O(n1332) );
  ND2CHD U1242 ( .I1(n1525), .I2(n1617), .O(n458) );
  AN2CHD U1243 ( .I1(n1524), .I2(n1523), .O(n1525) );
  ND2CHD U1244 ( .I1(rkey_next_17), .I2(n1584), .O(n1523) );
  ND2CHD U1245 ( .I1(n1852), .I2(rkey_next_33), .O(n1524) );
  AN2CHD U1246 ( .I1(n1679), .I2(n1678), .O(n1680) );
  AN2CHD U1247 ( .I1(n1674), .I2(n1673), .O(n1675) );
  AN2CHD U1248 ( .I1(n1670), .I2(n1669), .O(n1671) );
  ND2CHD U1249 ( .I1(n1852), .I2(rkey_next_20), .O(n1670) );
  ND2CHD U1250 ( .I1(n1807), .I2(Kin_20), .O(n1669) );
  ND2CHD U1251 ( .I1(n1543), .I2(n1611), .O(n462) );
  AN2CHD U1252 ( .I1(n1542), .I2(n1541), .O(n1543) );
  ND2CHD U1253 ( .I1(rkey_next_20), .I2(n1584), .O(n1541) );
  ND2CHD U1254 ( .I1(n1852), .I2(rkey_next_36), .O(n1542) );
  ND2CHD U1255 ( .I1(n1508), .I2(n1507), .O(n463) );
  ND2CHD U1256 ( .I1(n1506), .I2(n1852), .O(n1508) );
  AN2CHD U1257 ( .I1(n1666), .I2(n1665), .O(n1667) );
  ND2CHD U1258 ( .I1(n1851), .I2(key_39), .O(n1666) );
  AN2CHD U1259 ( .I1(n1657), .I2(n1656), .O(n1658) );
  ND2CHD U1260 ( .I1(n1852), .I2(rkey_next_23), .O(n1657) );
  ND2CHD U1261 ( .I1(n1807), .I2(Kin_23), .O(n1656) );
  ND2CHD U1262 ( .I1(n1347), .I2(n1605), .O(n466) );
  AN2CHD U1263 ( .I1(n1346), .I2(n1345), .O(n1347) );
  ND2CHD U1264 ( .I1(rkey_next_23), .I2(n1584), .O(n1345) );
  ND2CHD U1265 ( .I1(n1852), .I2(rkey_next_39), .O(n1346) );
  AN2CHD U1266 ( .I1(n1650), .I2(n1649), .O(n1651) );
  AN2CHD U1267 ( .I1(n1645), .I2(n1644), .O(n1646) );
  AN2CHD U1268 ( .I1(n1641), .I2(n1640), .O(n1642) );
  ND2CHD U1269 ( .I1(n1852), .I2(rkey_next_26), .O(n1641) );
  ND2CHD U1270 ( .I1(n1807), .I2(Kin_26), .O(n1640) );
  ND2CHD U1271 ( .I1(n1516), .I2(n1599), .O(n470) );
  AN2CHD U1272 ( .I1(n1515), .I2(n1514), .O(n1516) );
  ND2CHD U1273 ( .I1(rkey_next_26), .I2(n1584), .O(n1514) );
  ND2CHD U1274 ( .I1(n1852), .I2(rkey_next_42), .O(n1515) );
  AN2CHD U1275 ( .I1(n1634), .I2(n1633), .O(n1635) );
  ND2CHD U1276 ( .I1(n1851), .I2(key_45), .O(n1634) );
  AN2CHD U1277 ( .I1(n1625), .I2(n1624), .O(n1626) );
  ND2CHD U1278 ( .I1(n1852), .I2(rkey_next_29), .O(n1625) );
  ND2CHD U1279 ( .I1(n1540), .I2(n1593), .O(n474) );
  AN2CHD U1280 ( .I1(n1539), .I2(n1538), .O(n1540) );
  ND2CHD U1281 ( .I1(rkey_next_29), .I2(n1584), .O(n1538) );
  ND2CHD U1282 ( .I1(n1852), .I2(rkey_next_45), .O(n1539) );
  ND2CHD U1283 ( .I1(n1510), .I2(n1509), .O(n476) );
  ND2CHD U1284 ( .I1(n1852), .I2(rkey_next_16), .O(n1510) );
  ND2CHD U1285 ( .I1(n1546), .I2(n1619), .O(n477) );
  AN2CHD U1286 ( .I1(n1545), .I2(n1544), .O(n1546) );
  ND2CHD U1287 ( .I1(rkey_next_16), .I2(n1584), .O(n1544) );
  ND2CHD U1288 ( .I1(n1852), .I2(rkey_next_32), .O(n1545) );
  AN2CHD U1289 ( .I1(n1549), .I2(n1587), .O(n1550) );
  ND2CHD U1290 ( .I1(rkey_next_32), .I2(n1584), .O(n1549) );
  INVDHD U1291 ( .I(n869), .O(n824) );
  OR2EHD U1292 ( .I1(n764), .I2(n766), .O(n620) );
  AN2CHD U1293 ( .I1(n942), .I2(n941), .O(n623) );
  INVDHD U1294 ( .I(n797), .O(n1164) );
  ND2DHD U1295 ( .I1(n800), .I2(n799), .O(n797) );
  AN2CHD U1296 ( .I1(n1110), .I2(n782), .O(n624) );
  INVKHD U1297 ( .I(n631), .O(n718) );
  AN2HHD U1298 ( .I1(n819), .I2(n946), .O(n820) );
  INVGHD U1299 ( .I(n792), .O(n1156) );
  XNR3EHD U1300 ( .I1(n1242), .I2(n627), .I3(n1099), .O(n1128) );
  XNR3EHD U1301 ( .I1(n929), .I2(n928), .I3(n962), .O(n930) );
  OA22EHD U1302 ( .A1(n1285), .A2(n699), .B1(n1287), .B2(_keyexpantion_N26 ),.O(n1286) );
  XNR2KHD U1303 ( .I1(n1174), .I2(n1173), .O(n699) );
  OAI12CHD U1304 ( .B1(n1226), .B2(n1225), .A1(n628), .O(n629) );
  INVGHD U1305 ( .I(n1276), .O(n628) );
  XOR2HHD U1306 ( .I1(n956), .I2(n927), .O(n772) );
  XOR2HHD U1307 ( .I1(n1110), .I2(n636), .O(n927) );
  NR2GHD U1308 ( .I1(n869), .I2(n822), .O(n819) );
  INVGHD U1309 ( .I(n1058), .O(n709) );
  XNR2KHD U1310 ( .I1(n615), .I2(n629), .O(n677) );
  ND2KHD U1311 ( .I1(n630), .I2(n682), .O(n721) );
  ND3EHD U1312 ( .I1(n814), .I2(n812), .I3(n813), .O(n630) );
  INVGHD U1313 ( .I(n1057), .O(n708) );
  INVGHD U1314 ( .I(n1109), .O(n666) );
  INVHHD U1315 ( .I(n1287), .O(n631) );
  ND2KHD U1316 ( .I1(n1168), .I2(n1169), .O(n1183) );
  AN2HHD U1317 ( .I1(n840), .I2(n820), .O(n841) );
  INVLHD U1318 ( .I(n1329), .O(n935) );
  XNR3EHD U1319 ( .I1(n1021), .I2(n1029), .I3(n1031), .O(n1058) );
  NR2GHD U1320 ( .I1(n791), .I2(n808), .O(n807) );
  INVCKGHD U1321 ( .I(n1219), .O(n1220) );
  XNR2HHD U1322 ( .I1(n1189), .I2(n1199), .O(n1197) );
  INVDHD U1323 ( .I(n1291), .O(n725) );
  OAI22CHD U1324 ( .A1(n1060), .A2(n633), .B1(n644), .B2(n1054), .O(n1086) );
  ND3EHD U1325 ( .I1(n648), .I2(n647), .I3(n646), .O(n633) );
  XOR2HHD U1326 ( .I1(n1060), .I2(n633), .O(n643) );
  INVGHD U1327 ( .I(n634), .O(n1229) );
  ND2HHD U1328 ( .I1(n635), .I2(n1177), .O(n634) );
  ND2HHD U1329 ( .I1(n635), .I2(n752), .O(n684) );
  ND2HHD U1330 ( .I1(n1176), .I2(n635), .O(n1184) );
  ND2KHD U1331 ( .I1(n1170), .I2(n1171), .O(n635) );
  XNR2HHD U1332 ( .I1(n957), .I2(n959), .O(n956) );
  XOR2HHD U1333 ( .I1(n952), .I2(n1143), .O(n636) );
  XOR2HHD U1334 ( .I1(n1563), .I2(n773), .O(n1143) );
  ND2HHD U1335 ( .I1(n640), .I2(n639), .O(n1287) );
  ND3EHD U1336 ( .I1(n658), .I2(n1183), .I3(n1184), .O(n639) );
  ND2HHD U1337 ( .I1(n642), .I2(n641), .O(n640) );
  INVDHD U1338 ( .I(n1184), .O(n641) );
  ND2HHD U1339 ( .I1(n721), .I2(n1177), .O(n658) );
  ND2HHD U1340 ( .I1(n643), .I2(n722), .O(n776) );
  OAI22CHD U1341 ( .A1(n1086), .A2(n1085), .B1(n722), .B2(n643), .O(n707) );
  ND2DHD U1342 ( .I1(n1086), .I2(n1085), .O(n809) );
  MAOI1CHD U1343 ( .A1(n1052), .A2(n645), .B1(n1040), .B2(n1047), .O(n644) );
  ND3CHD U1344 ( .I1(n1053), .I2(n1078), .I3(n1054), .O(n646) );
  ND3EHD U1345 ( .I1(n645), .I2(n1052), .I3(n1051), .O(n647) );
  ND2DHD U1346 ( .I1(n697), .I2(n696), .O(n648) );
  XNR2HHD U1347 ( .I1(n1041), .I2(n649), .O(n1060) );
  XOR2HHD U1348 ( .I1(n1042), .I2(n1043), .O(n649) );
  XOR2HHD U1349 ( .I1(n626), .I2(n1547), .O(n1296) );
  ND2HHD U1350 ( .I1(n654), .I2(n650), .O(n1547) );
  ND3EHD U1351 ( .I1(n653), .I2(n652), .I3(n651), .O(n650) );
  ND2HHD U1352 ( .I1(n729), .I2(n1293), .O(n651) );
  ND2HHD U1353 ( .I1(n731), .I2(n730), .O(n653) );
  ND2HHD U1354 ( .I1(n656), .I2(n655), .O(n654) );
  NR2GHD U1355 ( .I1(n726), .I2(n723), .O(n655) );
  OAI12CHD U1356 ( .B1(n732), .B2(n677), .A1(n676), .O(n656) );
  ND2HHD U1357 ( .I1(n1059), .I2(n657), .O(n705) );
  XOR2HHD U1358 ( .I1(n1159), .I2(n1160), .O(n657) );
  NR2BHD U1359 ( .I1(n1175), .I2(n658), .O(n1182) );
  ND2HHD U1360 ( .I1(n1040), .I2(n1047), .O(n1052) );
  OA12HHD U1361 ( .B1(n661), .B2(n660), .A1(n659), .O(n1040) );
  ND2HHD U1362 ( .I1(n1089), .I2(n704), .O(n659) );
  NR2GHD U1363 ( .I1(n1045), .I2(n1089), .O(n661) );
  OAI12CHD U1364 ( .B1(n1056), .B2(n1055), .A1(n815), .O(n1057) );
  XOR2HHD U1365 ( .I1(n1020), .I2(n662), .O(n1055) );
  XOR2HHD U1366 ( .I1(n1016), .I2(n1017), .O(n662) );
  XOR2HHD U1367 ( .I1(n1093), .I2(n1010), .O(n1016) );
  ND2HHD U1368 ( .I1(n664), .I2(n663), .O(n1003) );
  ND3EHD U1369 ( .I1(n622), .I2(n1002), .I3(n999), .O(n663) );
  ND2HHD U1370 ( .I1(n747), .I2(n1041), .O(n664) );
  NR2IHD U1371 ( .I1(n618), .I2(n667), .O(n1157) );
  XOR2HHD U1372 ( .I1(n1167), .I2(n668), .O(n1169) );
  ND2KHD U1373 ( .I1(n692), .I2(n688), .O(n668) );
  MUX2HHD U1374 ( .A(n672), .B(n671), .S(n996), .O(n669) );
  ND2HHD U1375 ( .I1(n985), .I2(n670), .O(n996) );
  ND3CHD U1376 ( .I1(n974), .I2(n973), .I3(rnd_16), .O(n670) );
  XOR2HHD U1377 ( .I1(n976), .I2(n1319), .O(n985) );
  ND2HHD U1378 ( .I1(n1136), .I2(n993), .O(n672) );
  MXL2CHD U1379 ( .A(n674), .B(n675), .S(n1136), .OB(n673) );
  INVLHD U1380 ( .I(n994), .O(n1136) );
  XNR2HHD U1381 ( .I1(n972), .I2(n971), .O(n994) );
  NR2CHD U1382 ( .I1(n675), .I2(n993), .O(n674) );
  INVCKGHD U1383 ( .I(n995), .O(n675) );
  INVCKIHD U1384 ( .I(n677), .O(n1283) );
  ND2DHD U1385 ( .I1(n1228), .I2(n677), .O(n676) );
  ND2HHD U1386 ( .I1(n677), .I2(n1286), .O(n730) );
  ND2HHD U1387 ( .I1(n679), .I2(n678), .O(n1202) );
  AO12CHD U1388 ( .B1(n974), .B2(n824), .A1(n1350), .O(n679) );
  ND2HHD U1389 ( .I1(n680), .I2(n1291), .O(n1282) );
  INVCKIHD U1390 ( .I(n1288), .O(n680) );
  AN2HHD U1391 ( .I1(n1285), .I2(_keyexpantion_N26 ), .O(n1288) );
  XNR2CHD U1392 ( .I1(n1254), .I2(n1115), .O(n1253) );
  XNR2HHD U1393 ( .I1(n1115), .I2(n1118), .O(n1163) );
  ND2HHD U1394 ( .I1(n1225), .I2(n683), .O(n1173) );
  ND2HHD U1395 ( .I1(n721), .I2(n1229), .O(n1225) );
  NR2GHD U1396 ( .I1(n811), .I2(n807), .O(n682) );
  ND2HHD U1397 ( .I1(n684), .I2(n1176), .O(n1222) );
  ND2HHD U1398 ( .I1(n695), .I2(n1172), .O(n1176) );
  ND2HHD U1399 ( .I1(n685), .I2(n1553), .O(n803) );
  ND2HHD U1400 ( .I1(n806), .I2(n805), .O(n685) );
  ND2HHD U1401 ( .I1(n686), .I2(n797), .O(n805) );
  ND2HHD U1402 ( .I1(n1160), .I2(n687), .O(n806) );
  ND2HHD U1403 ( .I1(n756), .I2(n759), .O(n1160) );
  MUX2HHD U1404 ( .A(n690), .B(n689), .S(n785), .O(n688) );
  OAI12CHD U1405 ( .B1(n1022), .B2(n893), .A1(n894), .O(n689) );
  ND2CHD U1406 ( .I1(n1022), .I2(n893), .O(n691) );
  MUX2HHD U1407 ( .A(n693), .B(n617), .S(n1024), .O(n692) );
  ND2CHD U1408 ( .I1(n785), .I2(n1022), .O(n693) );
  XNR2KHD U1409 ( .I1(n1138), .I2(n825), .O(n785) );
  XOR2HHD U1410 ( .I1(n720), .I2(n694), .O(n1073) );
  ND2HHD U1411 ( .I1(n974), .I2(n839), .O(n694) );
  INVGHD U1412 ( .I(n1170), .O(n695) );
  XOR2HHD U1413 ( .I1(n1158), .I2(n1157), .O(n1170) );
  ND2DHD U1414 ( .I1(n1051), .I2(n1053), .O(n696) );
  NR2GHD U1415 ( .I1(n988), .I2(n1000), .O(n1043) );
  ND2HHD U1416 ( .I1(n1001), .I2(n998), .O(n1042) );
  INVMHD U1417 ( .I(n699), .O(n1291) );
  OA22EHD U1418 ( .A1(n1227), .A2(n699), .B1(n1287), .B2(n1857), .O(n1228) );
  INVCHD U1419 ( .I(n1072), .O(n703) );
  INVGHD U1420 ( .I(n1089), .O(n1077) );
  INVCHD U1421 ( .I(n1090), .O(n704) );
  NR2EHD U1422 ( .I1(n707), .I2(n791), .O(n814) );
  ND2HHD U1423 ( .I1(n706), .I2(n705), .O(n791) );
  ND2HHD U1424 ( .I1(n709), .I2(n708), .O(n706) );
  XOR2HHD U1425 ( .I1(n1055), .I2(n1056), .O(n1085) );
  AN2HHD U1426 ( .I1(n741), .I2(n619), .O(n1059) );
  ND3EHD U1427 ( .I1(n714), .I2(n713), .I3(n710), .O(n734) );
  MXL2CHD U1428 ( .A(n1271), .B(n1275), .S(n1274), .OB(n713) );
  MAOI1CHD U1429 ( .A1(n1274), .A2(n1273), .B1(n1278), .B2(n1277), .O(n714) );
  INVCHD U1430 ( .I(n1234), .O(n1248) );
  OAI22CHD U1431 ( .A1(n1265), .A2(n1264), .B1(n715), .B2(n1263), .O(n1266) );
  XNR2HHD U1432 ( .I1(n717), .I2(n716), .O(n1264) );
  XNR2HHD U1433 ( .I1(n1249), .I2(n1234), .O(n716) );
  INVDHD U1434 ( .I(n1263), .O(n717) );
  AN2HHD U1435 ( .I1(n1287), .I2(_keyexpantion_N26 ), .O(n728) );
  XOR2EHD U1436 ( .I1(n1036), .I2(n1037), .O(n720) );
  NR2EHD U1437 ( .I1(rnd_4), .I2(rnd_3), .O(n969) );
  ND3CHD U1438 ( .I1(n721), .I2(n1272), .I3(n1230), .O(n1231) );
  XNR2HHD U1439 ( .I1(n1185), .I2(n721), .O(n1285) );
  NR2BHD U1440 ( .I1(n721), .I2(n1179), .O(n1180) );
  ND2HHD U1441 ( .I1(n736), .I2(n1084), .O(n722) );
  ND2HHD U1442 ( .I1(n725), .I2(n1279), .O(n724) );
  ND2HHD U1443 ( .I1(n734), .I2(n727), .O(n726) );
  ND3EHD U1444 ( .I1(n728), .I2(n1291), .I3(n1280), .O(n727) );
  ND2HHD U1445 ( .I1(n1290), .I2(n1289), .O(n729) );
  ND2HHD U1446 ( .I1(n1284), .I2(n1283), .O(n731) );
  OAI22CHD U1447 ( .A1(n1291), .A2(n1187), .B1(n1186), .B2(n718), .O(n732) );
  OAI12CHD U1448 ( .B1(n614), .B2(n798), .A1(n733), .O(n760) );
  XOR2HHD U1449 ( .I1(n1252), .I2(n1026), .O(n1021) );
  XOR2HHD U1450 ( .I1(n1095), .I2(n1114), .O(n1026) );
  XOR2HHD U1451 ( .I1(n1561), .I2(n794), .O(n1114) );
  ND2HHD U1452 ( .I1(n1214), .I2(n1190), .O(n1095) );
  INVCHD U1453 ( .I(n1280), .O(n735) );
  ND2DHD U1454 ( .I1(n1087), .I2(n1088), .O(n736) );
  XNR3EHD U1455 ( .I1(n1080), .I2(n1079), .I3(n1078), .O(n1088) );
  XOR2HHD U1456 ( .I1(n909), .I2(n737), .O(n771) );
  XOR2CHD U1457 ( .I1(n737), .I2(n870), .O(n897) );
  ND2HHD U1458 ( .I1(n974), .I2(n973), .O(n737) );
  ND2DHD U1459 ( .I1(n738), .I2(n1042), .O(n747) );
  INVGHD U1460 ( .I(n1043), .O(n738) );
  XOR2HHD U1461 ( .I1(n986), .I2(n771), .O(n1062) );
  ND2HHD U1462 ( .I1(n743), .I2(n742), .O(n1102) );
  ND2HHD U1463 ( .I1(n1119), .I2(n1096), .O(n743) );
  ND2HHD U1464 ( .I1(n744), .I2(n1211), .O(n1119) );
  ND2HHD U1465 ( .I1(n1144), .I2(rnd_28), .O(n744) );
  ND2CHD U1466 ( .I1(n968), .I2(n969), .O(n746) );
  INVCKGHD U1467 ( .I(n1183), .O(n752) );
  ND2HHD U1468 ( .I1(n803), .I2(n804), .O(n1168) );
  XNR3EHD U1469 ( .I1(n922), .I2(n921), .I3(n772), .O(n1158) );
  XNR2HHD U1470 ( .I1(n1027), .I2(n753), .O(n1161) );
  ND2HHD U1471 ( .I1(n1009), .I2(n1008), .O(n753) );
  ND2HHD U1472 ( .I1(n1291), .I2(n1292), .O(n1293) );
  ND2HHD U1473 ( .I1(n718), .I2(n1281), .O(n1292) );
  NR2GHD U1474 ( .I1(_keyexpantion_N26 ), .I2(n1285), .O(n1281) );
  XOR2HHD U1475 ( .I1(n1122), .I2(n1123), .O(n1126) );
  ND2DHD U1476 ( .I1(n1091), .I2(n755), .O(n1011) );
  ND2DHD U1477 ( .I1(n1093), .I2(n755), .O(n1094) );
  OAI12CHD U1478 ( .B1(n757), .B2(n798), .A1(n797), .O(n756) );
  ND2HHD U1479 ( .I1(n760), .I2(n1164), .O(n759) );
  ND2KHD U1480 ( .I1(n937), .I2(n796), .O(n869) );
  NR2IHD U1481 ( .I1(rnd_11), .I2(rnd_10), .O(n796) );
  NR2IHD U1482 ( .I1(rnd_13), .I2(rnd_12), .O(n937) );
  ND2HHD U1483 ( .I1(n766), .I2(n765), .O(n1091) );
  ND2HHD U1484 ( .I1(n1010), .I2(n1093), .O(n1012) );
  ND3EHD U1485 ( .I1(n620), .I2(n763), .I3(n761), .O(n1010) );
  ND2DHD U1486 ( .I1(n762), .I2(n982), .O(n761) );
  INVGHD U1487 ( .I(n982), .O(n764) );
  ND3EHD U1488 ( .I1(n940), .I2(n942), .I3(n625), .O(n765) );
  AO12HHD U1489 ( .B1(n623), .B2(n940), .A1(n767), .O(n766) );
  XOR2HHD U1490 ( .I1(n1107), .I2(n1108), .O(n1093) );
  ND2CHD U1491 ( .I1(n946), .I2(n945), .O(n1107) );
  ND2HHD U1492 ( .I1(n768), .I2(n864), .O(n801) );
  ND2HHD U1493 ( .I1(n768), .I2(n908), .O(n783) );
  XOR2HHD U1494 ( .I1(n1188), .I2(n1193), .O(n964) );
  XNR2HHD U1495 ( .I1(n1195), .I2(n769), .O(n1193) );
  XNR3EHD U1496 ( .I1(n1204), .I2(n1198), .I3(n770), .O(n769) );
  XOR2EHD U1497 ( .I1(n1190), .I2(n1205), .O(n770) );
  MAO222CHD U1498 ( .A1(n772), .B1(n962), .C1(n963), .O(n1188) );
  ND2HHD U1499 ( .I1(n1177), .I2(n1183), .O(n1185) );
  OR3HHD U1500 ( .I1(n779), .I2(n778), .I3(n792), .O(n812) );
  ND2HHD U1501 ( .I1(n776), .I2(n777), .O(n792) );
  ND2HHD U1502 ( .I1(n1152), .I2(n1151), .O(n777) );
  NR2CHD U1503 ( .I1(n1150), .I2(n1149), .O(n778) );
  XNR2HHD U1504 ( .I1(n1128), .I2(n1127), .O(n1150) );
  OAI22CHD U1505 ( .A1(n784), .A2(n624), .B1(n781), .B2(n1133), .O(n1122) );
  INVCHD U1506 ( .I(n1132), .O(n781) );
  ND2CHD U1507 ( .I1(n1111), .I2(n1109), .O(n782) );
  XNR2KHD U1508 ( .I1(rnd_27), .I2(n783), .O(n1110) );
  OAI22CHD U1509 ( .A1(n1112), .A2(n1132), .B1(n1111), .B2(n793), .O(n784) );
  XOR2HHD U1510 ( .I1(n914), .I2(n632), .O(n977) );
  INVGHD U1511 ( .I(n1054), .O(n1051) );
  XNR2KHD U1512 ( .I1(n1032), .I2(n1110), .O(n1054) );
  XOR2HHD U1513 ( .I1(n1130), .I2(n1135), .O(n1032) );
  XOR2HHD U1514 ( .I1(n1557), .I2(n916), .O(n1135) );
  XOR2HHD U1515 ( .I1(n793), .I2(n920), .O(n1130) );
  INVCHD U1516 ( .I(rnd_17), .O(n793) );
  XOR2HHD U1517 ( .I1(n795), .I2(n1107), .O(n1214) );
  INVCHD U1518 ( .I(rnd_13), .O(n795) );
  AN2CHD U1519 ( .I1(n796), .I2(n1557), .O(n945) );
  ND2HHD U1520 ( .I1(n917), .I2(n796), .O(n1315) );
  ND2CHD U1521 ( .I1(n946), .I2(n796), .O(n916) );
  XNR3EHD U1522 ( .I1(n1105), .I2(n1092), .I3(n970), .O(n1020) );
  ND2DHD U1523 ( .I1(n1066), .I2(n1025), .O(n799) );
  ND2DHD U1524 ( .I1(n1026), .I2(n1252), .O(n800) );
  XNR2KHD U1525 ( .I1(rnd_30), .I2(n801), .O(n1250) );
  NR2GHD U1526 ( .I1(n802), .I2(n910), .O(n840) );
  ND2HHD U1527 ( .I1(n936), .I2(n934), .O(n910) );
  NR2EHD U1528 ( .I1(rnd_21), .I2(rnd_20), .O(n936) );
  NR2EHD U1529 ( .I1(rnd_23), .I2(rnd_22), .O(n872) );
  ND3EHD U1530 ( .I1(n806), .I2(_keyexpantion_N27 ), .I3(n805), .O(n804) );
  ND2KHD U1531 ( .I1(n842), .I2(n933), .O(n975) );
  NR2IHD U1532 ( .I1(rnd_5), .I2(rnd_4), .O(n933) );
  NR2IHD U1533 ( .I1(rnd_3), .I2(rnd_2), .O(n842) );
  XNR3EHD U1534 ( .I1(n1035), .I2(n990), .I3(n1140), .O(n1078) );
  AN2HHD U1535 ( .I1(n810), .I2(n809), .O(n808) );
  ND2HHD U1536 ( .I1(n1155), .I2(n1156), .O(n813) );
  NR2EHD U1537 ( .I1(n1232), .I2(n1231), .O(n1273) );
  ND2CHD U1538 ( .I1(dat_next_8), .I2(dat_next_15), .O(n817) );
  XOR2CHD U1539 ( .I1(dat_next_14), .I2(Dout_0), .O(n816) );
  XNR2CHD U1540 ( .I1(n817), .I2(n816), .O(n818) );
  ND2KHD U1541 ( .I1(n840), .I2(n871), .O(n1033) );
  NR2IHD U1542 ( .I1(rnd_9), .I2(rnd_8), .O(n1306) );
  NR2IHD U1543 ( .I1(rnd_7), .I2(rnd_6), .O(n943) );
  NR2IHD U1544 ( .I1(n932), .I2(n975), .O(n946) );
  INVKHD U1545 ( .I(rnd_15), .O(n1559) );
  ND2KHD U1546 ( .I1(n1559), .I2(n1350), .O(n868) );
  ND2HHD U1547 ( .I1(n917), .I2(n1305), .O(n822) );
  INVGHD U1548 ( .I(n989), .O(n1138) );
  BUFNHD U1549 ( .I(n946), .O(n974) );
  XNR2KHD U1550 ( .I1(n1556), .I2(n974), .O(n1137) );
  ND2HHD U1551 ( .I1(n1137), .I2(n1038), .O(n912) );
  XOR2HHD U1552 ( .I1(n912), .I2(n1140), .O(n825) );
  INVDHD U1553 ( .I(n1038), .O(n827) );
  XNR2KHD U1554 ( .I1(n827), .I2(n826), .O(n1251) );
  NR2IHD U1555 ( .I1(n878), .I2(n869), .O(n834) );
  ND2DHD U1556 ( .I1(n917), .I2(n1560), .O(n830) );
  ND3CHD U1557 ( .I1(n834), .I2(n832), .I3(n829), .O(n838) );
  ND3CHD U1558 ( .I1(n832), .I2(n943), .I3(n831), .O(n833) );
  INVGHD U1559 ( .I(n834), .O(n835) );
  AN3HHD U1560 ( .I1(n838), .I2(n837), .I3(n836), .O(n1044) );
  INVGHD U1561 ( .I(n1044), .O(n890) );
  XNR2HHD U1562 ( .I1(n890), .I2(n1039), .O(n1244) );
  XNR2KHD U1563 ( .I1(n1251), .I2(n1244), .O(n1022) );
  XNR2KHD U1564 ( .I1(n1564), .I2(n841), .O(n1115) );
  ND3CHD U1565 ( .I1(n935), .I2(n853), .I3(n968), .O(n844) );
  XOR2HHD U1566 ( .I1(n935), .I2(rnd_9), .O(n845) );
  XOR2EHD U1567 ( .I1(n846), .I2(n845), .O(n1069) );
  INVCHD U1568 ( .I(n1069), .O(n847) );
  ND2DHD U1569 ( .I1(n848), .I2(n847), .O(n850) );
  ND2HHD U1570 ( .I1(n850), .I2(n849), .O(n1024) );
  ND3CHD U1571 ( .I1(n872), .I2(n851), .I3(n1564), .O(n852) );
  XOR2HHD U1572 ( .I1(rnd_4), .I2(n935), .O(n1215) );
  BUFGHD U1573 ( .I(n933), .O(n915) );
  XOR2CHD U1574 ( .I1(rnd_9), .I2(rnd_25), .O(n855) );
  OAI12CHD U1575 ( .B1(n879), .B2(n854), .A1(n855), .O(n859) );
  INVCHD U1576 ( .I(n855), .O(n857) );
  ND3CHD U1577 ( .I1(n857), .I2(n856), .I3(n915), .O(n858) );
  ND3CHD U1578 ( .I1(n859), .I2(n1215), .I3(n858), .O(n860) );
  XOR2HHD U1579 ( .I1(n877), .I2(n862), .O(n883) );
  NR2EHD U1580 ( .I1(rnd_26), .I2(rnd_27), .O(n1013) );
  NR2BHD U1581 ( .I1(rnd_28), .I2(rnd_29), .O(n863) );
  NR2EHD U1582 ( .I1(n874), .I2(n1033), .O(n864) );
  XOR2HHD U1583 ( .I1(n883), .I2(n1250), .O(n1023) );
  INVDHD U1584 ( .I(n1023), .O(n894) );
  NR2BHD U1585 ( .I1(rnd_10), .I2(rnd_7), .O(n865) );
  ND3CHD U1586 ( .I1(n872), .I2(n871), .I3(n1568), .O(n873) );
  OR3CHD U1587 ( .I1(n874), .I2(n910), .I3(n873), .O(n875) );
  NR2EHD U1588 ( .I1(n879), .I2(n878), .O(n880) );
  XNR2EHD U1589 ( .I1(n1555), .I2(n880), .O(n1240) );
  ND2HHD U1590 ( .I1(n1240), .I2(n1215), .O(n1071) );
  INVCHD U1591 ( .I(n1071), .O(n881) );
  INVDHD U1592 ( .I(n883), .O(n884) );
  INVDHD U1593 ( .I(n890), .O(n1045) );
  MAO222CHD U1594 ( .A1(n1022), .B1(n894), .C1(n893), .O(n895) );
  INVCHD U1595 ( .I(n897), .O(n900) );
  NR2EHD U1596 ( .I1(rnd_31), .I2(n898), .O(n987) );
  INVCHD U1597 ( .I(n987), .O(n899) );
  ND2HHD U1598 ( .I1(n999), .I2(n901), .O(n963) );
  XOR2HHD U1599 ( .I1(rnd_2), .I2(n963), .O(n922) );
  ND2HHD U1600 ( .I1(n907), .I2(n925), .O(n921) );
  NR2EHD U1601 ( .I1(rnd_26), .I2(n1033), .O(n908) );
  ND3EHD U1602 ( .I1(n935), .I2(n915), .I3(n914), .O(n971) );
  ND2CHD U1603 ( .I1(n937), .I2(n909), .O(n918) );
  ND2DHD U1604 ( .I1(n946), .I2(n919), .O(n920) );
  XNR3EHD U1605 ( .I1(n950), .I2(n1135), .I3(n666), .O(n957) );
  INVDHD U1606 ( .I(n1158), .O(n931) );
  INVGHD U1607 ( .I(n927), .O(n961) );
  XOR2HHD U1608 ( .I1(n963), .I2(n961), .O(n928) );
  OA22EHD U1609 ( .A1(n1157), .A2(n931), .B1(n930), .B2(rnd_2), .O(n965) );
  NR2EHD U1610 ( .I1(n932), .I2(n1315), .O(n942) );
  NR2EHD U1611 ( .I1(n1316), .I2(n975), .O(n944) );
  XOR2EHD U1612 ( .I1(n1144), .I2(n1210), .O(n1198) );
  INVCHD U1613 ( .I(n1013), .O(n947) );
  ND2HHD U1614 ( .I1(n955), .I2(n954), .O(n1204) );
  ND2HHD U1615 ( .I1(n967), .I2(n966), .O(n1223) );
  ND2HHD U1616 ( .I1(n1230), .I2(n1223), .O(n1174) );
  ND2HHD U1617 ( .I1(n997), .I2(n1136), .O(n980) );
  ND2HHD U1618 ( .I1(n1143), .I2(n994), .O(n978) );
  ND2HHD U1619 ( .I1(n978), .I2(n1131), .O(n979) );
  ND2HHD U1620 ( .I1(n980), .I2(n979), .O(n1017) );
  INVDHD U1621 ( .I(n1130), .O(n1109) );
  ND2HHD U1622 ( .I1(n1012), .I2(n1011), .O(n1027) );
  XOR2HHD U1623 ( .I1(n614), .I2(n1161), .O(n1031) );
  INVCHD U1624 ( .I(rnd_28), .O(n1567) );
  ND2CHD U1625 ( .I1(n1013), .I2(n1567), .O(n1014) );
  INVDHD U1626 ( .I(n1016), .O(n1019) );
  INVGHD U1627 ( .I(n1017), .O(n1018) );
  MAO222HHD U1628 ( .A1(n1020), .B1(n1019), .C1(n1018), .O(n1029) );
  XNR3EHD U1629 ( .I1(n1024), .I2(n1023), .I3(n1022), .O(n1159) );
  INVCHD U1630 ( .I(n1095), .O(n1025) );
  XOR2HHD U1631 ( .I1(n1028), .I2(n1029), .O(n1030) );
  OAI12CHD U1632 ( .B1(n1034), .B2(n1033), .A1(n1565), .O(n1035) );
  XNR2KHD U1633 ( .I1(_keyexpantion_N26 ), .I2(n1137), .O(n1089) );
  XOR2CHD U1634 ( .I1(rnd_5), .I2(rnd_15), .O(n1036) );
  NR2CHD U1635 ( .I1(n1046), .I2(n1045), .O(n1076) );
  OAI12CHD U1636 ( .B1(n1566), .B2(n1098), .A1(n1074), .O(n1080) );
  OAI12CHD U1637 ( .B1(n1077), .B2(n1076), .A1(n1075), .O(n1079) );
  INVCHD U1638 ( .I(n1082), .O(n1083) );
  ND2DHD U1639 ( .I1(n1081), .I2(n1083), .O(n1084) );
  XOR2HHD U1640 ( .I1(n1088), .I2(n1087), .O(n1152) );
  XNR3EHD U1641 ( .I1(n1090), .I2(n1250), .I3(n1089), .O(n1101) );
  AN2HHD U1642 ( .I1(n1095), .I2(n1094), .O(n1117) );
  NR2BHD U1643 ( .I1(n1117), .I2(n1118), .O(n1097) );
  XOR2HHD U1644 ( .I1(n1101), .I2(n1102), .O(n1127) );
  BUFIHD U1645 ( .I(n1114), .O(n1247) );
  XNR3EHD U1646 ( .I1(n1116), .I2(n1247), .I3(n1115), .O(n1123) );
  XNR3EHD U1647 ( .I1(n1121), .I2(n1120), .I3(n1119), .O(n1129) );
  ND2CHD U1648 ( .I1(n1124), .I2(n1123), .O(n1125) );
  INVCHD U1649 ( .I(n1149), .O(n1154) );
  OAI22CHD U1650 ( .A1(n1154), .A2(n1153), .B1(n1152), .B2(n1151), .O(n1155));
  INVDHD U1651 ( .I(n1171), .O(n1172) );
  MXL2CHD U1652 ( .A(n1177), .B(n1183), .S(n1184), .OB(n1181) );
  INVCHD U1653 ( .I(n1185), .O(n1178) );
  AN2EHD U1654 ( .I1(n1184), .I2(n1178), .O(n1179) );
  OA13EHD U1655 ( .B1(n1182), .B2(n1181), .B3(n1180), .A1(_keyexpantion_N26 ),.O(n1187) );
  INVDHD U1656 ( .I(n1281), .O(n1186) );
  INVCHD U1657 ( .I(n1188), .O(n1194) );
  INVCHD U1658 ( .I(n1198), .O(n1189) );
  XOR2HHD U1659 ( .I1(n1195), .I2(n1197), .O(n1192) );
  INVCHD U1660 ( .I(n1190), .O(n1191) );
  OA22EHD U1661 ( .A1(n1194), .A2(n1193), .B1(n1192), .B2(n1191), .O(n1219) );
  INVDHD U1662 ( .I(n1195), .O(n1196) );
  ND2HHD U1663 ( .I1(n1197), .I2(n1196), .O(n1201) );
  ND2DHD U1664 ( .I1(n1199), .I2(n1198), .O(n1200) );
  XNR2EHD U1665 ( .I1(n1247), .I2(n1245), .O(n1234) );
  ND2DHD U1666 ( .I1(n1205), .I2(n1204), .O(n1209) );
  ND2HHD U1667 ( .I1(n1209), .I2(n1208), .O(n1233) );
  XNR3EHD U1668 ( .I1(n1249), .I2(n1215), .I3(n1263), .O(n1216) );
  XOR2HHD U1669 ( .I1(n1235), .I2(n1236), .O(n1218) );
  ND2HHD U1670 ( .I1(n1219), .I2(n1218), .O(n1272) );
  INVDHD U1671 ( .I(n1218), .O(n1221) );
  ND2DHD U1672 ( .I1(n1221), .I2(n1220), .O(n1270) );
  ND2HHD U1673 ( .I1(n1222), .I2(n1230), .O(n1224) );
  ND2HHD U1674 ( .I1(n1224), .I2(n1223), .O(n1276) );
  INVCHD U1675 ( .I(n1230), .O(n1226) );
  ND2CHD U1676 ( .I1(n1285), .I2(n1857), .O(n1227) );
  INVDHD U1677 ( .I(n1229), .O(n1232) );
  OAI22CHD U1678 ( .A1(n1239), .A2(n1238), .B1(n1237), .B2(n1236), .O(n1269));
  ND2CHD U1679 ( .I1(n1202), .I2(n1240), .O(n1241) );
  XOR2EHD U1680 ( .I1(n1242), .I2(n1241), .O(n1243) );
  OAI22CHD U1681 ( .A1(n1249), .A2(n1248), .B1(n1247), .B2(n1246), .O(n1261));
  OAI22CHD U1682 ( .A1(n1257), .A2(n1256), .B1(n1255), .B2(n1254), .O(n1258));
  XNR2CHD U1683 ( .I1(n1259), .I2(n1258), .O(n1260) );
  XNR2EHD U1684 ( .I1(n1267), .I2(n1266), .O(n1268) );
  XOR2HHD U1685 ( .I1(n1269), .I2(n1268), .O(n1274) );
  INVDHD U1686 ( .I(n1276), .O(n1277) );
  INVGHD U1687 ( .I(n718), .O(n1279) );
  ND2HHD U1688 ( .I1(n1292), .I2(n1282), .O(n1284) );
  ND2DHD U1689 ( .I1(n1288), .I2(n718), .O(n1290) );
  ND2HHD U1690 ( .I1(n1296), .I2(n1572), .O(n1300) );
  ND2HHD U1691 ( .I1(n1300), .I2(n1299), .O(n500) );
  NR2BHD U1692 ( .I1(rnd_31), .I2(sel), .O(n1302) );
  ND2CHD U1693 ( .I1(n1302), .I2(n1301), .O(n1322) );
  NR2BHD U1694 ( .I1(rnd_28), .I2(_keyexpantion_N27 ), .O(n1303) );
  ND2CHD U1695 ( .I1(n1304), .I2(n1303), .O(n1321) );
  NR2BHD U1696 ( .I1(n1308), .I2(n1307), .O(n1314) );
  AN4CHD U1697 ( .I1(n1312), .I2(n1311), .I3(n1310), .I4(n1309), .O(n1313) );
  AN2CHD U1698 ( .I1(n1314), .I2(n1313), .O(n1318) );
  ND3CHD U1699 ( .I1(n1319), .I2(n1318), .I3(n1317), .O(n1320) );
  NR3BHD U1700 ( .I1(n1322), .I2(n1321), .I3(n1320), .O(n1323) );
  MAOI1CHD U1701 ( .A1(EN), .A2(n1323), .B1(BSY), .B2(EN), .O(n480) );
  OA22CHD U1702 ( .A1(n1584), .A2(sel), .B1(Dvld), .B2(EN), .O(n481) );
  INVCHD U1703 ( .I(n1573), .O(n1324) );
  ND2CHD U1704 ( .I1(_keyexpantion_N26 ), .I2(n1324), .O(n1326) );
  ND2CHD U1705 ( .I1(rnd_31), .I2(EN), .O(n1325) );
  AO12CHD U1706 ( .B1(Kvld), .B2(n1584), .A1(n1807), .O(n483) );
  AOI22BHD U1707 ( .A1(Kin_17), .A2(n1807), .B1(rkey_next_1), .B2(n1584),.O(n1331) );
  MXL2CHD U1708 ( .A(n1350), .B(n1559), .S(n1570), .OB(n596) );
  AOI22BHD U1709 ( .A1(Din_18), .A2(n1573), .B1(dat_next_2), .B2(n1571), .O(n1359) );
  INVCHD U1710 ( .I(rkey_next_37), .O(n1744) );
  INVCHD U1711 ( .I(rkey_next_2), .O(n1764) );
  AOI22BHD U1712 ( .A1(rkey_next_2), .A2(rkey_next_37), .B1(n1744), .B2(n1764), .O(n1412) );
  INVCHD U1713 ( .I(n1412), .O(n1352) );
  INVCHD U1714 ( .I(rkey_2), .O(n1769) );
  INVCHD U1715 ( .I(rkey_next_38), .O(n1825) );
  INVCHD U1716 ( .I(rkey_next_3), .O(n1842) );
  AOI22BHD U1717 ( .A1(rkey_next_3), .A2(rkey_next_38), .B1(n1825), .B2(n1842), .O(n1380) );
  MUX2CHD U1718 ( .A(rkey_2), .B(n1769), .S(n1380), .O(n1351) );
  XOR2CHD U1719 ( .I1(dat_next_0), .I2(Dout_2), .O(n1355) );
  ND2CHD U1720 ( .I1(dat_next_10), .I2(dat_next_1), .O(n1354) );
  ND2CHD U1721 ( .I1(n1354), .I2(n1355), .O(n1353) );
  OAI12CHD U1722 ( .B1(n1355), .B2(n1354), .A1(n1353), .O(n1357) );
  ND2CHD U1723 ( .I1(n1758), .I2(n1357), .O(n1356) );
  OAI112BHD U1724 ( .C1(n1758), .C2(n1357), .A1(n1572), .B1(n1356), .O(n1358));
  AOI22BHD U1725 ( .A1(Din_27), .A2(n1573), .B1(dat_next_11), .B2(n1571),.O(n1369) );
  INVCHD U1726 ( .I(rkey_next_46), .O(n1696) );
  INVCHD U1727 ( .I(rkey_next_11), .O(n1716) );
  AOI22BHD U1728 ( .A1(rkey_next_11), .A2(rkey_next_46), .B1(n1696), .B2(n1716), .O(n1400) );
  INVCHD U1729 ( .I(n1400), .O(n1361) );
  INVCHD U1730 ( .I(rkey_11), .O(n1721) );
  INVCHD U1731 ( .I(rkey_next_47), .O(n1776) );
  INVCHD U1732 ( .I(rkey_next_12), .O(n1796) );
  AOI22BHD U1733 ( .A1(rkey_next_12), .A2(rkey_next_47), .B1(n1776), .B2(n1796), .O(n1390) );
  MUX2CHD U1734 ( .A(rkey_11), .B(n1721), .S(n1390), .O(n1360) );
  INVCHD U1735 ( .I(dat_next_10), .O(n1365) );
  MAOI1CHD U1736 ( .A1(dat_next_9), .A2(Dout_11), .B1(Dout_11), .B2(dat_next_9), .O(n1364) );
  INVCHD U1737 ( .I(dat_next_3), .O(n1363) );
  OAI12CHD U1738 ( .B1(n1365), .B2(n1363), .A1(n1364), .O(n1362) );
  OAI13BHD U1739 ( .B1(n1365), .B2(n1364), .B3(n1363), .A1(n1362), .O(n1367));
  ND2CHD U1740 ( .I1(n1710), .I2(n1367), .O(n1366) );
  OAI112BHD U1741 ( .C1(n1710), .C2(n1367), .A1(n1572), .B1(n1366), .O(n1368));
  AOI22BHD U1742 ( .A1(Din_23), .A2(n1573), .B1(dat_next_7), .B2(n1571), .O(n1378) );
  INVCHD U1743 ( .I(rkey_next_42), .O(n1639) );
  INVCHD U1744 ( .I(rkey_next_7), .O(n1659) );
  AOI22BHD U1745 ( .A1(rkey_next_7), .A2(rkey_next_42), .B1(n1639), .B2(n1659), .O(n1433) );
  INVCHD U1746 ( .I(n1433), .O(n1371) );
  INVCHD U1747 ( .I(rkey_7), .O(n1664) );
  INVCHD U1748 ( .I(rkey_next_43), .O(n1712) );
  INVCHD U1749 ( .I(rkey_next_8), .O(n1732) );
  AOI22BHD U1750 ( .A1(rkey_next_8), .A2(rkey_next_43), .B1(n1712), .B2(n1732), .O(n1486) );
  MUX2CHD U1751 ( .A(rkey_7), .B(n1664), .S(n1486), .O(n1370) );
  INVCHD U1752 ( .I(dat_next_15), .O(n1374) );
  MAOI1CHD U1753 ( .A1(dat_next_5), .A2(Dout_7), .B1(Dout_7), .B2(dat_next_5), .O(n1373) );
  INVCHD U1754 ( .I(dat_next_6), .O(n1477) );
  OAI12CHD U1755 ( .B1(n1374), .B2(n1477), .A1(n1373), .O(n1372) );
  OAI13BHD U1756 ( .B1(n1374), .B2(n1373), .B3(n1477), .A1(n1372), .O(n1376));
  ND2CHD U1757 ( .I1(n1653), .I2(n1376), .O(n1375) );
  OAI112BHD U1758 ( .C1(n1653), .C2(n1376), .A1(n1572), .B1(n1375), .O(n1377));
  AOI22BHD U1759 ( .A1(Din_19), .A2(n1573), .B1(dat_next_3), .B2(n1571), .O(n1388) );
  INVCHD U1760 ( .I(n1380), .O(n1381) );
  INVCHD U1761 ( .I(rkey_3), .O(n1850) );
  INVCHD U1762 ( .I(rkey_next_39), .O(n1655) );
  INVCHD U1763 ( .I(rkey_next_4), .O(n1672) );
  AOI22BHD U1764 ( .A1(rkey_next_4), .A2(rkey_next_39), .B1(n1655), .B2(n1672), .O(n1464) );
  MUX2CHD U1765 ( .A(rkey_3), .B(n1850), .S(n1464), .O(n1379) );
  MAOI1CHD U1766 ( .A1(dat_next_1), .A2(Dout_3), .B1(Dout_3), .B2(dat_next_1), .O(n1384) );
  ND2CHD U1767 ( .I1(dat_next_11), .I2(dat_next_2), .O(n1383) );
  ND2CHD U1768 ( .I1(n1383), .I2(n1384), .O(n1382) );
  OAI12CHD U1769 ( .B1(n1384), .B2(n1383), .A1(n1382), .O(n1386) );
  ND2CHD U1770 ( .I1(n1511), .I2(n1386), .O(n1385) );
  OAI112BHD U1771 ( .C1(n1511), .C2(n1386), .A1(n1572), .B1(n1385), .O(n1387));
  AOI22BHD U1772 ( .A1(Din_28), .A2(n1573), .B1(dat_next_12), .B2(n1571),.O(n1399) );
  INVCHD U1773 ( .I(n1390), .O(n1391) );
  INVCHD U1774 ( .I(rkey_12), .O(n1801) );
  MUX2CHD U1775 ( .A(rkey_12), .B(n1801), .S(n1453), .O(n1389) );
  INVCHD U1776 ( .I(dat_next_11), .O(n1395) );
  MAOI1CHD U1777 ( .A1(dat_next_10), .A2(Dout_12), .B1(Dout_12), .B2(dat_next_10), .O(n1394) );
  INVCHD U1778 ( .I(dat_next_4), .O(n1393) );
  OAI12CHD U1779 ( .B1(n1395), .B2(n1393), .A1(n1394), .O(n1392) );
  OAI13BHD U1780 ( .B1(n1395), .B2(n1394), .B3(n1393), .A1(n1392), .O(n1397));
  ND2CHD U1781 ( .I1(n1790), .I2(n1397), .O(n1396) );
  OAI112BHD U1782 ( .C1(n1790), .C2(n1397), .A1(n1572), .B1(n1396), .O(n1398));
  AOI22BHD U1783 ( .A1(Din_26), .A2(n1573), .B1(dat_next_10), .B2(n1571),.O(n1410) );
  INVCHD U1784 ( .I(rkey_next_45), .O(n1623) );
  INVCHD U1785 ( .I(rkey_next_10), .O(n1643) );
  AOI22BHD U1786 ( .A1(rkey_next_10), .A2(rkey_next_45), .B1(n1623), .B2(n1643), .O(n1422) );
  INVCHD U1787 ( .I(n1422), .O(n1402) );
  INVCHD U1788 ( .I(rkey_10), .O(n1648) );
  MUX2CHD U1789 ( .A(rkey_10), .B(n1648), .S(n1400), .O(n1401) );
  INVCHD U1790 ( .I(dat_next_9), .O(n1406) );
  MAOI1CHD U1791 ( .A1(dat_next_8), .A2(Dout_10), .B1(Dout_10), .B2(dat_next_8), .O(n1405) );
  INVCHD U1792 ( .I(dat_next_2), .O(n1404) );
  OAI12CHD U1793 ( .B1(n1406), .B2(n1404), .A1(n1405), .O(n1403) );
  OAI13BHD U1794 ( .B1(n1406), .B2(n1405), .B3(n1404), .A1(n1403), .O(n1408));
  ND2CHD U1795 ( .I1(n1637), .I2(n1408), .O(n1407) );
  OAI112BHD U1796 ( .C1(n1637), .C2(n1408), .A1(n1572), .B1(n1407), .O(n1409));
  AOI22BHD U1797 ( .A1(Din_17), .A2(n1573), .B1(dat_next_1), .B2(n1571), .O(n1421) );
  INVCHD U1798 ( .I(n1411), .O(n1414) );
  INVCHD U1799 ( .I(rkey_1), .O(n1689) );
  MAOI1CHD U1800 ( .A1(dat_next_15), .A2(Dout_1), .B1(Dout_1), .B2(dat_next_15), .O(n1417) );
  ND2CHD U1801 ( .I1(dat_next_0), .I2(dat_next_9), .O(n1416) );
  ND2CHD U1802 ( .I1(n1416), .I2(n1417), .O(n1415) );
  OAI12CHD U1803 ( .B1(n1417), .B2(n1416), .A1(n1415), .O(n1419) );
  ND2CHD U1804 ( .I1(n1682), .I2(n1419), .O(n1418) );
  OAI112BHD U1805 ( .C1(n1682), .C2(n1419), .A1(n1572), .B1(n1418), .O(n1420));
  AOI22BHD U1806 ( .A1(Din_25), .A2(n1573), .B1(dat_next_9), .B2(n1571), .O(n1432) );
  INVCHD U1807 ( .I(rkey_next_44), .O(n1792) );
  INVCHD U1808 ( .I(rkey_next_9), .O(n1813) );
  AOI22BHD U1809 ( .A1(rkey_next_9), .A2(rkey_next_44), .B1(n1792), .B2(n1813), .O(n1484) );
  INVCHD U1810 ( .I(n1484), .O(n1424) );
  INVCHD U1811 ( .I(rkey_9), .O(n1818) );
  MUX2CHD U1812 ( .A(rkey_9), .B(n1818), .S(n1422), .O(n1423) );
  INVCHD U1813 ( .I(dat_next_8), .O(n1428) );
  MAOI1CHD U1814 ( .A1(dat_next_7), .A2(Dout_9), .B1(Dout_9), .B2(dat_next_7), .O(n1427) );
  INVCHD U1815 ( .I(dat_next_1), .O(n1426) );
  OAI12CHD U1816 ( .B1(n1428), .B2(n1426), .A1(n1427), .O(n1425) );
  OAI13BHD U1817 ( .B1(n1428), .B2(n1427), .B3(n1426), .A1(n1425), .O(n1430));
  ND2CHD U1818 ( .I1(n1806), .I2(n1430), .O(n1429) );
  OAI112BHD U1819 ( .C1(n1806), .C2(n1430), .A1(n1572), .B1(n1429), .O(n1431));
  AOI22BHD U1820 ( .A1(Din_22), .A2(n1573), .B1(dat_next_6), .B2(n1571), .O(n1441) );
  INVCHD U1821 ( .I(rkey_next_41), .O(n1809) );
  INVCHD U1822 ( .I(rkey_next_6), .O(n1829) );
  AOI22BHD U1823 ( .A1(rkey_next_6), .A2(rkey_next_41), .B1(n1809), .B2(n1829), .O(n1442) );
  INVCHD U1824 ( .I(n1442), .O(n1435) );
  INVCHD U1825 ( .I(rkey_6), .O(n1834) );
  MUX2CHD U1826 ( .A(rkey_6), .B(n1834), .S(n1433), .O(n1434) );
  INVCHD U1827 ( .I(dat_next_14), .O(n1501) );
  MAOI1CHD U1828 ( .A1(dat_next_4), .A2(Dout_6), .B1(Dout_6), .B2(dat_next_4), .O(n1437) );
  INVCHD U1829 ( .I(dat_next_5), .O(n1455) );
  OAI12CHD U1830 ( .B1(n1501), .B2(n1455), .A1(n1437), .O(n1436) );
  OAI13BHD U1831 ( .B1(n1501), .B2(n1437), .B3(n1455), .A1(n1436), .O(n1439));
  ND2CHD U1832 ( .I1(n1823), .I2(n1439), .O(n1438) );
  OAI112BHD U1833 ( .C1(n1823), .C2(n1439), .A1(n1572), .B1(n1438), .O(n1440));
  AOI22BHD U1834 ( .A1(Din_21), .A2(n1573), .B1(dat_next_5), .B2(n1571), .O(n1451) );
  INVCHD U1835 ( .I(rkey_next_40), .O(n1728) );
  INVCHD U1836 ( .I(rkey_next_5), .O(n1748) );
  AOI22BHD U1837 ( .A1(rkey_next_5), .A2(rkey_next_40), .B1(n1728), .B2(n1748), .O(n1462) );
  INVCHD U1838 ( .I(n1462), .O(n1444) );
  INVCHD U1839 ( .I(rkey_5), .O(n1753) );
  MUX2CHD U1840 ( .A(rkey_5), .B(n1753), .S(n1442), .O(n1443) );
  MAOI1CHD U1841 ( .A1(dat_next_3), .A2(Dout_5), .B1(Dout_5), .B2(dat_next_3), .O(n1447) );
  ND2CHD U1842 ( .I1(dat_next_13), .I2(dat_next_4), .O(n1446) );
  ND2CHD U1843 ( .I1(n1446), .I2(n1447), .O(n1445) );
  OAI12CHD U1844 ( .B1(n1447), .B2(n1446), .A1(n1445), .O(n1449) );
  ND2CHD U1845 ( .I1(n1742), .I2(n1449), .O(n1448) );
  OAI112BHD U1846 ( .C1(n1742), .C2(n1449), .A1(n1572), .B1(n1448), .O(n1450));
  AOI22BHD U1847 ( .A1(Din_29), .A2(n1573), .B1(dat_next_13), .B2(n1571),.O(n1461) );
  INVCHD U1848 ( .I(rkey_13), .O(n1632) );
  INVCHD U1849 ( .I(rkey_next_33), .O(n1684) );
  INVCHD U1850 ( .I(rkey_next_14), .O(n1700) );
  AOI22BHD U1851 ( .A1(rkey_next_14), .A2(rkey_next_33), .B1(n1684), .B2(n1700), .O(n1474) );
  INVCHD U1852 ( .I(dat_next_12), .O(n1457) );
  MAOI1CHD U1853 ( .A1(dat_next_11), .A2(Dout_13), .B1(Dout_13), .B2(dat_next_11), .O(n1456) );
  OAI12CHD U1854 ( .B1(n1457), .B2(n1455), .A1(n1456), .O(n1454) );
  OAI13BHD U1855 ( .B1(n1457), .B2(n1456), .B3(n1455), .A1(n1454), .O(n1459));
  ND2CHD U1856 ( .I1(n1621), .I2(n1459), .O(n1458) );
  OAI112BHD U1857 ( .C1(n1621), .C2(n1459), .A1(n1572), .B1(n1458), .O(n1460));
  AOI22BHD U1858 ( .A1(Din_20), .A2(n1573), .B1(dat_next_4), .B2(n1571), .O(n1472) );
  INVCHD U1859 ( .I(n1464), .O(n1465) );
  INVCHD U1860 ( .I(rkey_4), .O(n1677) );
  MUX2CHD U1861 ( .A(rkey_4), .B(n1677), .S(n1462), .O(n1463) );
  MAOI1CHD U1862 ( .A1(dat_next_2), .A2(Dout_4), .B1(Dout_4), .B2(dat_next_2), .O(n1468) );
  ND2CHD U1863 ( .I1(dat_next_12), .I2(dat_next_3), .O(n1467) );
  ND2CHD U1864 ( .I1(n1467), .I2(n1468), .O(n1466) );
  OAI12CHD U1865 ( .B1(n1468), .B2(n1467), .A1(n1466), .O(n1470) );
  ND2CHD U1866 ( .I1(n1506), .I2(n1470), .O(n1469) );
  OAI112BHD U1867 ( .C1(n1506), .C2(n1470), .A1(n1572), .B1(n1469), .O(n1471));
  AOI22BHD U1868 ( .A1(dat_next_14), .A2(n1571), .B1(n1573), .B2(Din_30),.O(n1483) );
  INVCHD U1869 ( .I(n1474), .O(n1475) );
  INVCHD U1870 ( .I(rkey_14), .O(n1705) );
  INVCHD U1871 ( .I(rkey_next_34), .O(n1760) );
  INVCHD U1872 ( .I(rkey_next_15), .O(n1780) );
  AOI22BHD U1873 ( .A1(rkey_next_15), .A2(rkey_next_34), .B1(n1760), .B2(n1780), .O(n1495) );
  MUX2CHD U1874 ( .A(rkey_14), .B(n1705), .S(n1495), .O(n1473) );
  INVCHD U1875 ( .I(dat_next_13), .O(n1479) );
  MAOI1CHD U1876 ( .A1(dat_next_12), .A2(Dout_14), .B1(Dout_14), .B2(dat_next_12), .O(n1478) );
  OAI12CHD U1877 ( .B1(n1479), .B2(n1477), .A1(n1478), .O(n1476) );
  OAI13BHD U1878 ( .B1(n1479), .B2(n1478), .B3(n1477), .A1(n1476), .O(n1481));
  ND2CHD U1879 ( .I1(n1694), .I2(n1481), .O(n1480) );
  OAI112BHD U1880 ( .C1(n1694), .C2(n1481), .A1(n1572), .B1(n1480), .O(n1482));
  AOI22BHD U1881 ( .A1(dat_next_8), .A2(n1571), .B1(n1573), .B2(Din_24), .O(n1494) );
  INVCHD U1882 ( .I(n1486), .O(n1487) );
  INVCHD U1883 ( .I(rkey_8), .O(n1737) );
  MUX2CHD U1884 ( .A(rkey_8), .B(n1737), .S(n1484), .O(n1485) );
  MAOI1CHD U1885 ( .A1(dat_next_6), .A2(Dout_8), .B1(Dout_8), .B2(dat_next_6), .O(n1490) );
  INVCHD U1886 ( .I(dat_next_0), .O(n1488) );
  INVCHD U1887 ( .I(dat_next_7), .O(n1499) );
  OR2CHD U1888 ( .I1(n1488), .I2(n1499), .O(n1489) );
  XNR2CHD U1889 ( .I1(n1490), .I2(n1489), .O(n1492) );
  ND2CHD U1890 ( .I1(n1726), .I2(n1492), .O(n1491) );
  OAI112BHD U1891 ( .C1(n1726), .C2(n1492), .A1(n1572), .B1(n1491), .O(n1493));
  AOI22BHD U1892 ( .A1(dat_next_15), .A2(n1571), .B1(n1573), .B2(Din_31),.O(n1505) );
  MAOI1CHD U1893 ( .A1(n1495), .A2(rkey_15), .B1(rkey_15), .B2(n1495), .O(n1496) );
  MAOI1CHD U1894 ( .A1(dat_next_13), .A2(Dout_15), .B1(Dout_15), .B2(dat_next_13), .O(n1500) );
  OAI12CHD U1895 ( .B1(n1501), .B2(n1499), .A1(n1500), .O(n1498) );
  OAI13BHD U1896 ( .B1(n1501), .B2(n1500), .B3(n1499), .A1(n1498), .O(n1503));
  ND2CHD U1897 ( .I1(n1774), .I2(n1503), .O(n1502) );
  OAI112BHD U1898 ( .C1(n1774), .C2(n1503), .A1(n1572), .B1(n1502), .O(n1504));
  AOI22BHD U1899 ( .A1(Kin_52), .A2(n1807), .B1(rkey_next_36), .B2(n1584),.O(n1507) );
  AOI22BHD U1900 ( .A1(Kin_16), .A2(n1807), .B1(rkey_next_0), .B2(n1584),.O(n1509) );
  AOI22BHD U1901 ( .A1(Kin_51), .A2(n1807), .B1(rkey_next_35), .B2(n1584),.O(n1512) );
  XNR2HHD U1902 ( .I1(n1548), .I2(n1547), .O(n1552) );
  OAI12CHD U1903 ( .B1(n1552), .B2(n1551), .A1(n1550), .O(n478) );
  MXL2CHD U1904 ( .A(n1857), .B(n1553), .S(n1570), .OB(n610) );
  MXL2CHD U1905 ( .A(n1553), .B(n1579), .S(n1570), .OB(n609) );
  MXL2CHD U1906 ( .A(n1554), .B(n1555), .S(n1570), .OB(n602) );
  MXL2CHD U1907 ( .A(n1555), .B(n1556), .S(n1570), .OB(n601) );
  MXL2CHD U1908 ( .A(n1556), .B(n1558), .S(n1570), .OB(n600) );
  MXL2CHD U1909 ( .A(n1558), .B(n1557), .S(n1570), .OB(n599) );
  MXL2CHD U1910 ( .A(n1559), .B(n909), .S(n1570), .OB(n595) );
  MXL2CHD U1911 ( .A(n788), .B(n1563), .S(n1570), .OB(n589) );
  MXL2CHD U1912 ( .A(n1564), .B(n1566), .S(n1570), .OB(n586) );
  MXL2CHD U1913 ( .A(n1566), .B(n1565), .S(n1570), .OB(n585) );
  MXL2CHD U1914 ( .A(n1567), .B(n1569), .S(n1570), .OB(n582) );
  MXL2CHD U1915 ( .A(n1569), .B(n1568), .S(n1570), .OB(n581) );
  MUX2CHD U1916 ( .A(sel), .B(rnd_31), .S(EN), .O(n482) );
  ND2CHD U1917 ( .I1(n1573), .I2(Din_0), .O(n1574) );
  ND3CHD U1918 ( .I1(n1576), .I2(n1575), .I3(n1574), .O(n516) );
  INVCHD U1919 ( .I(rkey_next_0), .O(n1582) );
  AOI22BHD U1920 ( .A1(n1845), .A2(key_48), .B1(n1851), .B2(key_32), .O(n1581) );
  AOI22BHD U1921 ( .A1(n1807), .A2(Kin_0), .B1(rkey_0), .B2(n1584), .O(n1580) );
  OAI112BHD U1922 ( .C1(n1551), .C2(n1582), .A1(n1581), .B1(n1580), .O(n1586));
  NR3BHD U1923 ( .I1(Krdy), .I2(n1857), .I3(n1584), .O(n1843) );
  AOI22BHD U1924 ( .A1(n1844), .A2(key_16), .B1(n1843), .B2(key_0), .O(n1585) );
  OR2B1CHD U1925 ( .I1(n1586), .B1(n1585), .O(n479) );
  INVCHD U1926 ( .I(key_48), .O(n1588) );
  OAI12CHD U1927 ( .B1(n1807), .B2(n1588), .A1(n1587), .O(n565) );
  INVCHD U1928 ( .I(key_47), .O(n1590) );
  OAI12CHD U1929 ( .B1(n1807), .B2(n1590), .A1(n1589), .O(n564) );
  INVCHD U1930 ( .I(key_46), .O(n1592) );
  OAI12CHD U1931 ( .B1(n1807), .B2(n1592), .A1(n1591), .O(n563) );
  INVCHD U1932 ( .I(key_45), .O(n1594) );
  OAI12CHD U1933 ( .B1(n1807), .B2(n1594), .A1(n1593), .O(n562) );
  INVCHD U1934 ( .I(key_44), .O(n1596) );
  OAI12CHD U1935 ( .B1(n1807), .B2(n1596), .A1(n1595), .O(n561) );
  INVCHD U1936 ( .I(key_43), .O(n1598) );
  OAI12CHD U1937 ( .B1(n1807), .B2(n1598), .A1(n1597), .O(n560) );
  INVCHD U1938 ( .I(key_42), .O(n1600) );
  OAI12CHD U1939 ( .B1(n1807), .B2(n1600), .A1(n1599), .O(n559) );
  INVCHD U1940 ( .I(key_41), .O(n1602) );
  OAI12CHD U1941 ( .B1(n1807), .B2(n1602), .A1(n1601), .O(n558) );
  INVCHD U1942 ( .I(key_40), .O(n1604) );
  OAI12CHD U1943 ( .B1(n1807), .B2(n1604), .A1(n1603), .O(n557) );
  INVCHD U1944 ( .I(key_39), .O(n1606) );
  OAI12CHD U1945 ( .B1(n1807), .B2(n1606), .A1(n1605), .O(n556) );
  INVCHD U1946 ( .I(key_38), .O(n1608) );
  OAI12CHD U1947 ( .B1(n1807), .B2(n1608), .A1(n1607), .O(n555) );
  INVCHD U1948 ( .I(key_37), .O(n1610) );
  OAI12CHD U1949 ( .B1(n1807), .B2(n1610), .A1(n1609), .O(n554) );
  INVCHD U1950 ( .I(key_36), .O(n1612) );
  OAI12CHD U1951 ( .B1(n1807), .B2(n1612), .A1(n1611), .O(n553) );
  INVCHD U1952 ( .I(key_35), .O(n1614) );
  OAI12CHD U1953 ( .B1(n1807), .B2(n1614), .A1(n1613), .O(n552) );
  INVCHD U1954 ( .I(key_34), .O(n1616) );
  OAI12CHD U1955 ( .B1(n1807), .B2(n1616), .A1(n1615), .O(n551) );
  INVCHD U1956 ( .I(key_33), .O(n1618) );
  OAI12CHD U1957 ( .B1(n1807), .B2(n1618), .A1(n1617), .O(n550) );
  INVCHD U1958 ( .I(key_32), .O(n1620) );
  OAI12CHD U1959 ( .B1(n1807), .B2(n1620), .A1(n1619), .O(n549) );
  AOI22BHD U1960 ( .A1(n1807), .A2(Kin_61), .B1(n1621), .B2(n1852), .O(n1622));
  OAI12CHD U1961 ( .B1(EN), .B2(n1623), .A1(n1622), .O(n475) );
  INVCHD U1962 ( .I(rkey_next_13), .O(n1627) );
  OAI12CHD U1963 ( .B1(EN), .B2(n1627), .A1(n1626), .O(n473) );
  AOI22BHD U1964 ( .A1(n1844), .A2(key_29), .B1(n1843), .B2(key_13), .O(n1631) );
  OAI112BHD U1965 ( .C1(EN), .C2(n1632), .A1(n1631), .B1(n1630), .O(n1636) );
  OR2B1CHD U1966 ( .I1(n1636), .B1(n1635), .O(n472) );
  AOI22BHD U1967 ( .A1(n1807), .A2(Kin_58), .B1(n1637), .B2(n1852), .O(n1638));
  OAI12CHD U1968 ( .B1(EN), .B2(n1639), .A1(n1638), .O(n471) );
  OAI12CHD U1969 ( .B1(EN), .B2(n1643), .A1(n1642), .O(n469) );
  AOI22BHD U1970 ( .A1(n1844), .A2(key_26), .B1(n1843), .B2(key_10), .O(n1647) );
  ND2CHD U1971 ( .I1(n1807), .I2(Kin_10), .O(n1644) );
  OAI112BHD U1972 ( .C1(EN), .C2(n1648), .A1(n1647), .B1(n1646), .O(n1652) );
  OR2B1CHD U1973 ( .I1(n1652), .B1(n1651), .O(n468) );
  AOI22BHD U1974 ( .A1(n1807), .A2(Kin_55), .B1(n1653), .B2(n1852), .O(n1654));
  OAI12CHD U1975 ( .B1(EN), .B2(n1655), .A1(n1654), .O(n467) );
  OAI12CHD U1976 ( .B1(EN), .B2(n1659), .A1(n1658), .O(n465) );
  AOI22BHD U1977 ( .A1(n1844), .A2(key_23), .B1(n1843), .B2(key_7), .O(n1663) );
  OAI112BHD U1978 ( .C1(EN), .C2(n1664), .A1(n1663), .B1(n1662), .O(n1668) );
  OR2B1CHD U1979 ( .I1(n1668), .B1(n1667), .O(n464) );
  OAI12CHD U1980 ( .B1(EN), .B2(n1672), .A1(n1671), .O(n461) );
  AOI22BHD U1981 ( .A1(n1844), .A2(key_20), .B1(n1843), .B2(key_4), .O(n1676) );
  ND2CHD U1982 ( .I1(n1807), .I2(Kin_4), .O(n1673) );
  OAI112BHD U1983 ( .C1(EN), .C2(n1677), .A1(n1676), .B1(n1675), .O(n1681) );
  OR2B1CHD U1984 ( .I1(n1681), .B1(n1680), .O(n460) );
  AOI22BHD U1985 ( .A1(n1807), .A2(Kin_49), .B1(n1682), .B2(n1852), .O(n1683));
  OAI12CHD U1986 ( .B1(EN), .B2(n1684), .A1(n1683), .O(n459) );
  AOI22BHD U1987 ( .A1(n1844), .A2(key_17), .B1(n1843), .B2(key_1), .O(n1688) );
  ND2CHD U1988 ( .I1(n1807), .I2(Kin_1), .O(n1685) );
  OAI112BHD U1989 ( .C1(EN), .C2(n1689), .A1(n1688), .B1(n1687), .O(n1693) );
  OR2B1CHD U1990 ( .I1(n1693), .B1(n1692), .O(n456) );
  AOI22BHD U1991 ( .A1(n1807), .A2(Kin_62), .B1(n1694), .B2(n1852), .O(n1695));
  OAI12CHD U1992 ( .B1(EN), .B2(n1696), .A1(n1695), .O(n455) );
  OAI12CHD U1993 ( .B1(EN), .B2(n1700), .A1(n1699), .O(n453) );
  AOI22BHD U1994 ( .A1(n1844), .A2(key_30), .B1(n1843), .B2(key_14), .O(n1704) );
  ND2CHD U1995 ( .I1(n1807), .I2(Kin_14), .O(n1701) );
  OAI112BHD U1996 ( .C1(EN), .C2(n1705), .A1(n1704), .B1(n1703), .O(n1709) );
  OR2B1CHD U1997 ( .I1(n1709), .B1(n1708), .O(n452) );
  AOI22BHD U1998 ( .A1(n1807), .A2(Kin_59), .B1(n1710), .B2(n1852), .O(n1711));
  OAI12CHD U1999 ( .B1(EN), .B2(n1712), .A1(n1711), .O(n451) );
  OAI12CHD U2000 ( .B1(EN), .B2(n1716), .A1(n1715), .O(n449) );
  AOI22BHD U2001 ( .A1(n1844), .A2(key_27), .B1(n1843), .B2(key_11), .O(n1720) );
  ND2CHD U2002 ( .I1(n1807), .I2(Kin_11), .O(n1717) );
  OAI112BHD U2003 ( .C1(EN), .C2(n1721), .A1(n1720), .B1(n1719), .O(n1725) );
  OR2B1CHD U2004 ( .I1(n1725), .B1(n1724), .O(n448) );
  AOI22BHD U2005 ( .A1(n1807), .A2(Kin_56), .B1(n1726), .B2(n1852), .O(n1727));
  OAI12CHD U2006 ( .B1(EN), .B2(n1728), .A1(n1727), .O(n447) );
  OAI12CHD U2007 ( .B1(EN), .B2(n1732), .A1(n1731), .O(n445) );
  AOI22BHD U2008 ( .A1(n1844), .A2(key_24), .B1(n1843), .B2(key_8), .O(n1736) );
  OAI112BHD U2009 ( .C1(EN), .C2(n1737), .A1(n1736), .B1(n1735), .O(n1741) );
  OR2B1CHD U2010 ( .I1(n1741), .B1(n1740), .O(n444) );
  AOI22BHD U2011 ( .A1(n1807), .A2(Kin_53), .B1(n1742), .B2(n1852), .O(n1743));
  OAI12CHD U2012 ( .B1(EN), .B2(n1744), .A1(n1743), .O(n443) );
  OAI12CHD U2013 ( .B1(EN), .B2(n1748), .A1(n1747), .O(n441) );
  AOI22BHD U2014 ( .A1(n1844), .A2(key_21), .B1(n1843), .B2(key_5), .O(n1752) );
  ND2CHD U2015 ( .I1(n1807), .I2(Kin_5), .O(n1749) );
  OAI112BHD U2016 ( .C1(EN), .C2(n1753), .A1(n1752), .B1(n1751), .O(n1757) );
  OR2B1CHD U2017 ( .I1(n1757), .B1(n1756), .O(n440) );
  AOI22BHD U2018 ( .A1(n1807), .A2(Kin_50), .B1(n1758), .B2(n1852), .O(n1759));
  OAI12CHD U2019 ( .B1(EN), .B2(n1760), .A1(n1759), .O(n439) );
  OAI12CHD U2020 ( .B1(EN), .B2(n1764), .A1(n1763), .O(n437) );
  AOI22BHD U2021 ( .A1(n1844), .A2(key_18), .B1(n1843), .B2(key_2), .O(n1768) );
  OAI112BHD U2022 ( .C1(EN), .C2(n1769), .A1(n1768), .B1(n1767), .O(n1773) );
  OR2B1CHD U2023 ( .I1(n1773), .B1(n1772), .O(n436) );
  AOI22BHD U2024 ( .A1(n1807), .A2(Kin_63), .B1(n1774), .B2(n1852), .O(n1775));
  OAI12CHD U2025 ( .B1(EN), .B2(n1776), .A1(n1775), .O(n435) );
  OAI12CHD U2026 ( .B1(EN), .B2(n1780), .A1(n1779), .O(n433) );
  INVCHD U2027 ( .I(rkey_15), .O(n1785) );
  AOI22BHD U2028 ( .A1(n1844), .A2(key_31), .B1(n1843), .B2(key_15), .O(n1784) );
  OAI112BHD U2029 ( .C1(EN), .C2(n1785), .A1(n1784), .B1(n1783), .O(n1789) );
  OR2B1CHD U2030 ( .I1(n1789), .B1(n1788), .O(n432) );
  AOI22BHD U2031 ( .A1(n1807), .A2(Kin_60), .B1(n1790), .B2(n1852), .O(n1791));
  OAI12CHD U2032 ( .B1(EN), .B2(n1792), .A1(n1791), .O(n431) );
  OAI12CHD U2033 ( .B1(EN), .B2(n1796), .A1(n1795), .O(n429) );
  AOI22BHD U2034 ( .A1(n1844), .A2(key_28), .B1(n1843), .B2(key_12), .O(n1800) );
  OAI112BHD U2035 ( .C1(EN), .C2(n1801), .A1(n1800), .B1(n1799), .O(n1805) );
  OR2B1CHD U2036 ( .I1(n1805), .B1(n1804), .O(n428) );
  AOI22BHD U2037 ( .A1(n1807), .A2(Kin_57), .B1(n1806), .B2(n1852), .O(n1808));
  OAI12CHD U2038 ( .B1(EN), .B2(n1809), .A1(n1808), .O(n427) );
  OAI12CHD U2039 ( .B1(EN), .B2(n1813), .A1(n1812), .O(n425) );
  AOI22BHD U2040 ( .A1(n1844), .A2(key_25), .B1(n1843), .B2(key_9), .O(n1817) );
  ND2CHD U2041 ( .I1(n1807), .I2(Kin_9), .O(n1814) );
  OAI112BHD U2042 ( .C1(EN), .C2(n1818), .A1(n1817), .B1(n1816), .O(n1822) );
  OR2B1CHD U2043 ( .I1(n1822), .B1(n1821), .O(n424) );
  AOI22BHD U2044 ( .A1(n1807), .A2(Kin_54), .B1(n1823), .B2(n1852), .O(n1824));
  OAI12CHD U2045 ( .B1(EN), .B2(n1825), .A1(n1824), .O(n423) );
  OAI12CHD U2046 ( .B1(EN), .B2(n1829), .A1(n1828), .O(n421) );
  AOI22BHD U2047 ( .A1(n1844), .A2(key_22), .B1(n1843), .B2(key_6), .O(n1833) );
  ND2CHD U2048 ( .I1(n1807), .I2(Kin_6), .O(n1830) );
  OAI112BHD U2049 ( .C1(EN), .C2(n1834), .A1(n1833), .B1(n1832), .O(n1838) );
  OR2B1CHD U2050 ( .I1(n1838), .B1(n1837), .O(n420) );
  OAI12CHD U2051 ( .B1(EN), .B2(n1842), .A1(n1841), .O(n417) );
  AOI22BHD U2052 ( .A1(n1844), .A2(key_19), .B1(n1843), .B2(key_3), .O(n1849) );
  OAI112BHD U2053 ( .C1(EN), .C2(n1850), .A1(n1849), .B1(n1848), .O(n1856) );
  OR2B1CHD U2054 ( .I1(n1856), .B1(n1855), .O(n416) );
  BUFCHD U2055 ( .I1(Dout_31), .O(dat_next_15) );
  BUFCHD U2056 ( .I1(Dout_30), .O(dat_next_14) );
  BUFCHD U2057 ( .I1(Dout_29), .O(dat_next_13) );
  BUFCHD U2058 ( .I1(Dout_28), .O(dat_next_12) );
  BUFCHD U2059 ( .I1(Dout_27), .O(dat_next_11) );
  BUFCHD U2060 ( .I1(Dout_26), .O(dat_next_10) );
  BUFCHD U2061 ( .I1(Dout_25), .O(dat_next_9) );
  BUFCHD U2062 ( .I1(Dout_24), .O(dat_next_8) );
  BUFCHD U2063 ( .I1(Dout_23), .O(dat_next_7) );
  BUFCHD U2064 ( .I1(Dout_22), .O(dat_next_6) );
  BUFCHD U2065 ( .I1(Dout_21), .O(dat_next_5) );
  BUFCHD U2066 ( .I1(Dout_20), .O(dat_next_4) );
  BUFCHD U2067 ( .I1(Dout_19), .O(dat_next_3) );
  BUFCHD U2068 ( .I1(Dout_18), .O(dat_next_2) );
  BUFCHD U2069 ( .I1(Dout_17), .O(dat_next_1) );
  BUFCHD U2070 ( .I1(Dout_16), .O(dat_next_0) );
endmodule


