module CLEFIA ( 
CLK, 
SRST, 
MODE_0,
MODE_1,
ENCDEC, 
KEYSET, 
DATASET, 
KEY_0,
KEY_1,
KEY_2,
KEY_3,
KEY_4,
KEY_5,
KEY_6,
KEY_7,
KEY_8,
KEY_9,
KEY_10,
KEY_11,
KEY_12,
KEY_13,
KEY_14,
KEY_15,
KEY_16,
KEY_17,
KEY_18,
KEY_19,
KEY_20,
KEY_21,
KEY_22,
KEY_23,
KEY_24,
KEY_25,
KEY_26,
KEY_27,
KEY_28,
KEY_29,
KEY_30,
KEY_31,
KEY_32,
KEY_33,
KEY_34,
KEY_35,
KEY_36,
KEY_37,
KEY_38,
KEY_39,
KEY_40,
KEY_41,
KEY_42,
KEY_43,
KEY_44,
KEY_45,
KEY_46,
KEY_47,
KEY_48,
KEY_49,
KEY_50,
KEY_51,
KEY_52,
KEY_53,
KEY_54,
KEY_55,
KEY_56,
KEY_57,
KEY_58,
KEY_59,
KEY_60,
KEY_61,
KEY_62,
KEY_63,
KEY_64,
KEY_65,
KEY_66,
KEY_67,
KEY_68,
KEY_69,
KEY_70,
KEY_71,
KEY_72,
KEY_73,
KEY_74,
KEY_75,
KEY_76,
KEY_77,
KEY_78,
KEY_79,
KEY_80,
KEY_81,
KEY_82,
KEY_83,
KEY_84,
KEY_85,
KEY_86,
KEY_87,
KEY_88,
KEY_89,
KEY_90,
KEY_91,
KEY_92,
KEY_93,
KEY_94,
KEY_95,
KEY_96,
KEY_97,
KEY_98,
KEY_99,
KEY_100,
KEY_101,
KEY_102,
KEY_103,
KEY_104,
KEY_105,
KEY_106,
KEY_107,
KEY_108,
KEY_109,
KEY_110,
KEY_111,
KEY_112,
KEY_113,
KEY_114,
KEY_115,
KEY_116,
KEY_117,
KEY_118,
KEY_119,
KEY_120,
KEY_121,
KEY_122,
KEY_123,
KEY_124,
KEY_125,
KEY_126,
KEY_127,
KEY_128,
KEY_129,
KEY_130,
KEY_131,
KEY_132,
KEY_133,
KEY_134,
KEY_135,
KEY_136,
KEY_137,
KEY_138,
KEY_139,
KEY_140,
KEY_141,
KEY_142,
KEY_143,
KEY_144,
KEY_145,
KEY_146,
KEY_147,
KEY_148,
KEY_149,
KEY_150,
KEY_151,
KEY_152,
KEY_153,
KEY_154,
KEY_155,
KEY_156,
KEY_157,
KEY_158,
KEY_159,
KEY_160,
KEY_161,
KEY_162,
KEY_163,
KEY_164,
KEY_165,
KEY_166,
KEY_167,
KEY_168,
KEY_169,
KEY_170,
KEY_171,
KEY_172,
KEY_173,
KEY_174,
KEY_175,
KEY_176,
KEY_177,
KEY_178,
KEY_179,
KEY_180,
KEY_181,
KEY_182,
KEY_183,
KEY_184,
KEY_185,
KEY_186,
KEY_187,
KEY_188,
KEY_189,
KEY_190,
KEY_191,
KEY_192,
KEY_193,
KEY_194,
KEY_195,
KEY_196,
KEY_197,
KEY_198,
KEY_199,
KEY_200,
KEY_201,
KEY_202,
KEY_203,
KEY_204,
KEY_205,
KEY_206,
KEY_207,
KEY_208,
KEY_209,
KEY_210,
KEY_211,
KEY_212,
KEY_213,
KEY_214,
KEY_215,
KEY_216,
KEY_217,
KEY_218,
KEY_219,
KEY_220,
KEY_221,
KEY_222,
KEY_223,
KEY_224,
KEY_225,
KEY_226,
KEY_227,
KEY_228,
KEY_229,
KEY_230,
KEY_231,
KEY_232,
KEY_233,
KEY_234,
KEY_235,
KEY_236,
KEY_237,
KEY_238,
KEY_239,
KEY_240,
KEY_241,
KEY_242,
KEY_243,
KEY_244,
KEY_245,
KEY_246,
KEY_247,
KEY_248,
KEY_249,
KEY_250,
KEY_251,
KEY_252,
KEY_253,
KEY_254,
KEY_255,
DIN_0,
DIN_1,
DIN_2,
DIN_3,
DIN_4,
DIN_5,
DIN_6,
DIN_7,
DIN_8,
DIN_9,
DIN_10,
DIN_11,
DIN_12,
DIN_13,
DIN_14,
DIN_15,
DIN_16,
DIN_17,
DIN_18,
DIN_19,
DIN_20,
DIN_21,
DIN_22,
DIN_23,
DIN_24,
DIN_25,
DIN_26,
DIN_27,
DIN_28,
DIN_29,
DIN_30,
DIN_31,
DIN_32,
DIN_33,
DIN_34,
DIN_35,
DIN_36,
DIN_37,
DIN_38,
DIN_39,
DIN_40,
DIN_41,
DIN_42,
DIN_43,
DIN_44,
DIN_45,
DIN_46,
DIN_47,
DIN_48,
DIN_49,
DIN_50,
DIN_51,
DIN_52,
DIN_53,
DIN_54,
DIN_55,
DIN_56,
DIN_57,
DIN_58,
DIN_59,
DIN_60,
DIN_61,
DIN_62,
DIN_63,
DIN_64,
DIN_65,
DIN_66,
DIN_67,
DIN_68,
DIN_69,
DIN_70,
DIN_71,
DIN_72,
DIN_73,
DIN_74,
DIN_75,
DIN_76,
DIN_77,
DIN_78,
DIN_79,
DIN_80,
DIN_81,
DIN_82,
DIN_83,
DIN_84,
DIN_85,
DIN_86,
DIN_87,
DIN_88,
DIN_89,
DIN_90,
DIN_91,
DIN_92,
DIN_93,
DIN_94,
DIN_95,
DIN_96,
DIN_97,
DIN_98,
DIN_99,
DIN_100,
DIN_101,
DIN_102,
DIN_103,
DIN_104,
DIN_105,
DIN_106,
DIN_107,
DIN_108,
DIN_109,
DIN_110,
DIN_111,
DIN_112,
DIN_113,
DIN_114,
DIN_115,
DIN_116,
DIN_117,
DIN_118,
DIN_119,
DIN_120,
DIN_121,
DIN_122,
DIN_123,
DIN_124,
DIN_125,
DIN_126,
DIN_127,
BSY, 
DVLD, 
DOUT_0,
DOUT_1,
DOUT_2,
DOUT_3,
DOUT_4,
DOUT_5,
DOUT_6,
DOUT_7,
DOUT_8,
DOUT_9,
DOUT_10,
DOUT_11,
DOUT_12,
DOUT_13,
DOUT_14,
DOUT_15,
DOUT_16,
DOUT_17,
DOUT_18,
DOUT_19,
DOUT_20,
DOUT_21,
DOUT_22,
DOUT_23,
DOUT_24,
DOUT_25,
DOUT_26,
DOUT_27,
DOUT_28,
DOUT_29,
DOUT_30,
DOUT_31,
DOUT_32,
DOUT_33,
DOUT_34,
DOUT_35,
DOUT_36,
DOUT_37,
DOUT_38,
DOUT_39,
DOUT_40,
DOUT_41,
DOUT_42,
DOUT_43,
DOUT_44,
DOUT_45,
DOUT_46,
DOUT_47,
DOUT_48,
DOUT_49,
DOUT_50,
DOUT_51,
DOUT_52,
DOUT_53,
DOUT_54,
DOUT_55,
DOUT_56,
DOUT_57,
DOUT_58,
DOUT_59,
DOUT_60,
DOUT_61,
DOUT_62,
DOUT_63,
DOUT_64,
DOUT_65,
DOUT_66,
DOUT_67,
DOUT_68,
DOUT_69,
DOUT_70,
DOUT_71,
DOUT_72,
DOUT_73,
DOUT_74,
DOUT_75,
DOUT_76,
DOUT_77,
DOUT_78,
DOUT_79,
DOUT_80,
DOUT_81,
DOUT_82,
DOUT_83,
DOUT_84,
DOUT_85,
DOUT_86,
DOUT_87,
DOUT_88,
DOUT_89,
DOUT_90,
DOUT_91,
DOUT_92,
DOUT_93,
DOUT_94,
DOUT_95,
DOUT_96,
DOUT_97,
DOUT_98,
DOUT_99,
DOUT_100,
DOUT_101,
DOUT_102,
DOUT_103,
DOUT_104,
DOUT_105,
DOUT_106,
DOUT_107,
DOUT_108,
DOUT_109,
DOUT_110,
DOUT_111,
DOUT_112,
DOUT_113,
DOUT_114,
DOUT_115,
DOUT_116,
DOUT_117,
DOUT_118,
DOUT_119,
DOUT_120,
DOUT_121,
DOUT_122,
DOUT_123,
DOUT_124,
DOUT_125,
DOUT_126,
DOUT_127
);
//Start PIs
input MODE_0;
input MODE_1;
input KEY_0;
input KEY_1;
input KEY_2;
input KEY_3;
input KEY_4;
input KEY_5;
input KEY_6;
input KEY_7;
input KEY_8;
input KEY_9;
input KEY_10;
input KEY_11;
input KEY_12;
input KEY_13;
input KEY_14;
input KEY_15;
input KEY_16;
input KEY_17;
input KEY_18;
input KEY_19;
input KEY_20;
input KEY_21;
input KEY_22;
input KEY_23;
input KEY_24;
input KEY_25;
input KEY_26;
input KEY_27;
input KEY_28;
input KEY_29;
input KEY_30;
input KEY_31;
input KEY_32;
input KEY_33;
input KEY_34;
input KEY_35;
input KEY_36;
input KEY_37;
input KEY_38;
input KEY_39;
input KEY_40;
input KEY_41;
input KEY_42;
input KEY_43;
input KEY_44;
input KEY_45;
input KEY_46;
input KEY_47;
input KEY_48;
input KEY_49;
input KEY_50;
input KEY_51;
input KEY_52;
input KEY_53;
input KEY_54;
input KEY_55;
input KEY_56;
input KEY_57;
input KEY_58;
input KEY_59;
input KEY_60;
input KEY_61;
input KEY_62;
input KEY_63;
input KEY_64;
input KEY_65;
input KEY_66;
input KEY_67;
input KEY_68;
input KEY_69;
input KEY_70;
input KEY_71;
input KEY_72;
input KEY_73;
input KEY_74;
input KEY_75;
input KEY_76;
input KEY_77;
input KEY_78;
input KEY_79;
input KEY_80;
input KEY_81;
input KEY_82;
input KEY_83;
input KEY_84;
input KEY_85;
input KEY_86;
input KEY_87;
input KEY_88;
input KEY_89;
input KEY_90;
input KEY_91;
input KEY_92;
input KEY_93;
input KEY_94;
input KEY_95;
input KEY_96;
input KEY_97;
input KEY_98;
input KEY_99;
input KEY_100;
input KEY_101;
input KEY_102;
input KEY_103;
input KEY_104;
input KEY_105;
input KEY_106;
input KEY_107;
input KEY_108;
input KEY_109;
input KEY_110;
input KEY_111;
input KEY_112;
input KEY_113;
input KEY_114;
input KEY_115;
input KEY_116;
input KEY_117;
input KEY_118;
input KEY_119;
input KEY_120;
input KEY_121;
input KEY_122;
input KEY_123;
input KEY_124;
input KEY_125;
input KEY_126;
input KEY_127;
input KEY_128;
input KEY_129;
input KEY_130;
input KEY_131;
input KEY_132;
input KEY_133;
input KEY_134;
input KEY_135;
input KEY_136;
input KEY_137;
input KEY_138;
input KEY_139;
input KEY_140;
input KEY_141;
input KEY_142;
input KEY_143;
input KEY_144;
input KEY_145;
input KEY_146;
input KEY_147;
input KEY_148;
input KEY_149;
input KEY_150;
input KEY_151;
input KEY_152;
input KEY_153;
input KEY_154;
input KEY_155;
input KEY_156;
input KEY_157;
input KEY_158;
input KEY_159;
input KEY_160;
input KEY_161;
input KEY_162;
input KEY_163;
input KEY_164;
input KEY_165;
input KEY_166;
input KEY_167;
input KEY_168;
input KEY_169;
input KEY_170;
input KEY_171;
input KEY_172;
input KEY_173;
input KEY_174;
input KEY_175;
input KEY_176;
input KEY_177;
input KEY_178;
input KEY_179;
input KEY_180;
input KEY_181;
input KEY_182;
input KEY_183;
input KEY_184;
input KEY_185;
input KEY_186;
input KEY_187;
input KEY_188;
input KEY_189;
input KEY_190;
input KEY_191;
input KEY_192;
input KEY_193;
input KEY_194;
input KEY_195;
input KEY_196;
input KEY_197;
input KEY_198;
input KEY_199;
input KEY_200;
input KEY_201;
input KEY_202;
input KEY_203;
input KEY_204;
input KEY_205;
input KEY_206;
input KEY_207;
input KEY_208;
input KEY_209;
input KEY_210;
input KEY_211;
input KEY_212;
input KEY_213;
input KEY_214;
input KEY_215;
input KEY_216;
input KEY_217;
input KEY_218;
input KEY_219;
input KEY_220;
input KEY_221;
input KEY_222;
input KEY_223;
input KEY_224;
input KEY_225;
input KEY_226;
input KEY_227;
input KEY_228;
input KEY_229;
input KEY_230;
input KEY_231;
input KEY_232;
input KEY_233;
input KEY_234;
input KEY_235;
input KEY_236;
input KEY_237;
input KEY_238;
input KEY_239;
input KEY_240;
input KEY_241;
input KEY_242;
input KEY_243;
input KEY_244;
input KEY_245;
input KEY_246;
input KEY_247;
input KEY_248;
input KEY_249;
input KEY_250;
input KEY_251;
input KEY_252;
input KEY_253;
input KEY_254;
input KEY_255;
input DIN_0;
input DIN_1;
input DIN_2;
input DIN_3;
input DIN_4;
input DIN_5;
input DIN_6;
input DIN_7;
input DIN_8;
input DIN_9;
input DIN_10;
input DIN_11;
input DIN_12;
input DIN_13;
input DIN_14;
input DIN_15;
input DIN_16;
input DIN_17;
input DIN_18;
input DIN_19;
input DIN_20;
input DIN_21;
input DIN_22;
input DIN_23;
input DIN_24;
input DIN_25;
input DIN_26;
input DIN_27;
input DIN_28;
input DIN_29;
input DIN_30;
input DIN_31;
input DIN_32;
input DIN_33;
input DIN_34;
input DIN_35;
input DIN_36;
input DIN_37;
input DIN_38;
input DIN_39;
input DIN_40;
input DIN_41;
input DIN_42;
input DIN_43;
input DIN_44;
input DIN_45;
input DIN_46;
input DIN_47;
input DIN_48;
input DIN_49;
input DIN_50;
input DIN_51;
input DIN_52;
input DIN_53;
input DIN_54;
input DIN_55;
input DIN_56;
input DIN_57;
input DIN_58;
input DIN_59;
input DIN_60;
input DIN_61;
input DIN_62;
input DIN_63;
input DIN_64;
input DIN_65;
input DIN_66;
input DIN_67;
input DIN_68;
input DIN_69;
input DIN_70;
input DIN_71;
input DIN_72;
input DIN_73;
input DIN_74;
input DIN_75;
input DIN_76;
input DIN_77;
input DIN_78;
input DIN_79;
input DIN_80;
input DIN_81;
input DIN_82;
input DIN_83;
input DIN_84;
input DIN_85;
input DIN_86;
input DIN_87;
input DIN_88;
input DIN_89;
input DIN_90;
input DIN_91;
input DIN_92;
input DIN_93;
input DIN_94;
input DIN_95;
input DIN_96;
input DIN_97;
input DIN_98;
input DIN_99;
input DIN_100;
input DIN_101;
input DIN_102;
input DIN_103;
input DIN_104;
input DIN_105;
input DIN_106;
input DIN_107;
input DIN_108;
input DIN_109;
input DIN_110;
input DIN_111;
input DIN_112;
input DIN_113;
input DIN_114;
input DIN_115;
input DIN_116;
input DIN_117;
input DIN_118;
input DIN_119;
input DIN_120;
input DIN_121;
input DIN_122;
input DIN_123;
input DIN_124;
input DIN_125;
input DIN_126;
input DIN_127;
input CLK;
input SRST;
input ENCDEC;
input KEYSET;
input DATASET;
//Start POs
output DOUT_0;
output DOUT_1;
output DOUT_2;
output DOUT_3;
output DOUT_4;
output DOUT_5;
output DOUT_6;
output DOUT_7;
output DOUT_8;
output DOUT_9;
output DOUT_10;
output DOUT_11;
output DOUT_12;
output DOUT_13;
output DOUT_14;
output DOUT_15;
output DOUT_16;
output DOUT_17;
output DOUT_18;
output DOUT_19;
output DOUT_20;
output DOUT_21;
output DOUT_22;
output DOUT_23;
output DOUT_24;
output DOUT_25;
output DOUT_26;
output DOUT_27;
output DOUT_28;
output DOUT_29;
output DOUT_30;
output DOUT_31;
output DOUT_32;
output DOUT_33;
output DOUT_34;
output DOUT_35;
output DOUT_36;
output DOUT_37;
output DOUT_38;
output DOUT_39;
output DOUT_40;
output DOUT_41;
output DOUT_42;
output DOUT_43;
output DOUT_44;
output DOUT_45;
output DOUT_46;
output DOUT_47;
output DOUT_48;
output DOUT_49;
output DOUT_50;
output DOUT_51;
output DOUT_52;
output DOUT_53;
output DOUT_54;
output DOUT_55;
output DOUT_56;
output DOUT_57;
output DOUT_58;
output DOUT_59;
output DOUT_60;
output DOUT_61;
output DOUT_62;
output DOUT_63;
output DOUT_64;
output DOUT_65;
output DOUT_66;
output DOUT_67;
output DOUT_68;
output DOUT_69;
output DOUT_70;
output DOUT_71;
output DOUT_72;
output DOUT_73;
output DOUT_74;
output DOUT_75;
output DOUT_76;
output DOUT_77;
output DOUT_78;
output DOUT_79;
output DOUT_80;
output DOUT_81;
output DOUT_82;
output DOUT_83;
output DOUT_84;
output DOUT_85;
output DOUT_86;
output DOUT_87;
output DOUT_88;
output DOUT_89;
output DOUT_90;
output DOUT_91;
output DOUT_92;
output DOUT_93;
output DOUT_94;
output DOUT_95;
output DOUT_96;
output DOUT_97;
output DOUT_98;
output DOUT_99;
output DOUT_100;
output DOUT_101;
output DOUT_102;
output DOUT_103;
output DOUT_104;
output DOUT_105;
output DOUT_106;
output DOUT_107;
output DOUT_108;
output DOUT_109;
output DOUT_110;
output DOUT_111;
output DOUT_112;
output DOUT_113;
output DOUT_114;
output DOUT_115;
output DOUT_116;
output DOUT_117;
output DOUT_118;
output DOUT_119;
output DOUT_120;
output DOUT_121;
output DOUT_122;
output DOUT_123;
output DOUT_124;
output DOUT_125;
output DOUT_126;
output DOUT_127;
output BSY;
output DVLD;
//Start wires
wire _i_CLEFIA128_CON_T_xi_2;
wire _i_CLEFIA128_CON_T_reg_4;
wire n6095;
wire n6096;
wire n6097;
wire n6098;
wire n6099;
wire n6100;
wire n6101;
wire n6102;
wire n6103;
wire n6104;
wire n6105;
wire n6106;
wire n6107;
wire n6108;
wire n6109;
wire n6110;
wire n6111;
wire n6112;
wire n6113;
wire n6114;
wire n6115;
wire n6116;
wire n6117;
wire n6118;
wire n6119;
wire n6120;
wire n6121;
wire n6122;
wire n6123;
wire n6124;
wire n6125;
wire n6126;
wire n6127;
wire n6128;
wire n6129;
wire n6130;
wire n6131;
wire n6132;
wire n6133;
wire n6134;
wire n6135;
wire n6136;
wire n6137;
wire n6138;
wire n6139;
wire n6140;
wire n6141;
wire n6142;
wire n6143;
wire n6144;
wire n6145;
wire n6146;
wire n6147;
wire n6148;
wire n6149;
wire n6150;
wire n6151;
wire n6152;
wire n6153;
wire n6154;
wire n6155;
wire n6156;
wire n6157;
wire n6158;
wire n6159;
wire n6160;
wire n6161;
wire n6162;
wire n6163;
wire n6164;
wire n6165;
wire n6166;
wire n6167;
wire n6168;
wire n6169;
wire n6170;
wire n6171;
wire n6172;
wire n6173;
wire n6174;
wire n6175;
wire n6176;
wire n6177;
wire n6178;
wire n6179;
wire n6180;
wire n6181;
wire n6182;
wire n6183;
wire n6184;
wire n6185;
wire n6186;
wire n6187;
wire n6188;
wire n6189;
wire n6190;
wire n6191;
wire n6192;
wire n6193;
wire n6194;
wire n6195;
wire n6196;
wire n6197;
wire n6198;
wire n6199;
wire n6200;
wire n6201;
wire n6202;
wire n6203;
wire n6204;
wire n6205;
wire n6206;
wire n6207;
wire n6208;
wire n6209;
wire n6210;
wire n6211;
wire n6212;
wire n6213;
wire n6214;
wire n6215;
wire n6216;
wire n6217;
wire n6218;
wire n6219;
wire n6220;
wire n6221;
wire n6222;
wire n6223;
wire n6224;
wire n6225;
wire n6226;
wire n6227;
wire n6228;
wire n6229;
wire n6230;
wire n6231;
wire n6232;
wire n6233;
wire n6234;
wire n6235;
wire n6236;
wire n6237;
wire n6238;
wire n6239;
wire n6240;
wire n6241;
wire n6242;
wire n6243;
wire n6244;
wire n6245;
wire n6246;
wire n6247;
wire n6248;
wire n6249;
wire n6250;
wire n6251;
wire n6252;
wire n6253;
wire n6254;
wire n6255;
wire n6256;
wire n6257;
wire n6258;
wire n6259;
wire n6260;
wire n6261;
wire n6262;
wire n6263;
wire n6264;
wire n6265;
wire n6266;
wire n6267;
wire n6268;
wire n6269;
wire n6270;
wire n6271;
wire n6272;
wire n6273;
wire n6274;
wire n6275;
wire n6276;
wire n6277;
wire n6278;
wire n6279;
wire n6280;
wire n6281;
wire n6282;
wire n6283;
wire n6284;
wire n6285;
wire n6286;
wire n6287;
wire n6288;
wire n6289;
wire n6290;
wire n6291;
wire n6292;
wire n6293;
wire n6294;
wire n6295;
wire n6296;
wire n6297;
wire n6298;
wire n6299;
wire n6300;
wire n6301;
wire n6302;
wire n6303;
wire n6304;
wire n6305;
wire n6306;
wire n6307;
wire n6308;
wire n6309;
wire n6310;
wire n6311;
wire n6312;
wire n6313;
wire n6314;
wire n6315;
wire n6316;
wire n6317;
wire n6318;
wire n6319;
wire n6320;
wire n6321;
wire n6322;
wire n6323;
wire n6324;
wire n6325;
wire n6326;
wire n6327;
wire n6328;
wire n6329;
wire n6330;
wire n6331;
wire n6332;
wire n6333;
wire n6334;
wire n6335;
wire n6336;
wire n6337;
wire n6338;
wire n6339;
wire n6340;
wire n6341;
wire n6342;
wire n6343;
wire n6344;
wire n6345;
wire n6346;
wire n6347;
wire n6348;
wire n6349;
wire n6350;
wire n6351;
wire n6352;
wire n6353;
wire n6354;
wire n6355;
wire n6356;
wire n6357;
wire n6358;
wire n6359;
wire n6360;
wire n6361;
wire n6362;
wire n6363;
wire n6364;
wire n6365;
wire n6366;
wire n6367;
wire n6368;
wire n6370;
wire n6371;
wire n6372;
wire n6373;
wire n6374;
wire n6375;
wire n6376;
wire n6377;
wire n6378;
wire n6379;
wire n6380;
wire n6381;
wire n6382;
wire n6383;
wire n6384;
wire n6385;
wire n6386;
wire n6387;
wire n6388;
wire n6389;
wire n6390;
wire n6391;
wire n6392;
wire n6393;
wire n6394;
wire n6395;
wire n6396;
wire n6397;
wire n6398;
wire n6399;
wire n6400;
wire n6401;
wire n6402;
wire n6403;
wire n6404;
wire n6405;
wire n6406;
wire n6407;
wire n6408;
wire n6409;
wire n6410;
wire n6411;
wire n6412;
wire n6413;
wire n6414;
wire n6415;
wire n6416;
wire n6417;
wire n6418;
wire n6419;
wire n6420;
wire n6421;
wire n6422;
wire n6423;
wire n6424;
wire n6425;
wire n6426;
wire n6427;
wire n6428;
wire n6429;
wire n6430;
wire n6431;
wire n6432;
wire n6433;
wire n6434;
wire n6435;
wire n6436;
wire n6437;
wire n6438;
wire n6439;
wire n6440;
wire n6441;
wire n6442;
wire n6443;
wire n6444;
wire n6445;
wire n6446;
wire n6447;
wire n6448;
wire n6449;
wire n6450;
wire n6451;
wire n6452;
wire n6453;
wire n6454;
wire n6455;
wire n6456;
wire n6457;
wire n6458;
wire n6459;
wire n6460;
wire n6461;
wire n6462;
wire n6463;
wire n6464;
wire n6465;
wire n6466;
wire n6467;
wire n6468;
wire n6469;
wire n6470;
wire n6471;
wire n6472;
wire n6473;
wire n6474;
wire n6475;
wire n6476;
wire n6477;
wire n6478;
wire n6479;
wire n6480;
wire n6481;
wire n6482;
wire n6483;
wire n6484;
wire n6485;
wire n6486;
wire n6487;
wire n6488;
wire n6489;
wire n6490;
wire n6491;
wire n6492;
wire n6493;
wire n6494;
wire n6495;
wire n6496;
wire n6497;
wire n6498;
wire n6499;
wire n6500;
wire n6501;
wire n6502;
wire n6503;
wire n6504;
wire n6505;
wire n6506;
wire n6507;
wire n6508;
wire n6509;
wire n6510;
wire n6511;
wire n6512;
wire n6513;
wire n6514;
wire n6515;
wire n6516;
wire n6517;
wire n6518;
wire n6519;
wire n6520;
wire n6521;
wire n6522;
wire n6523;
wire n6524;
wire n6525;
wire n6526;
wire n6527;
wire n6528;
wire n6529;
wire n6530;
wire n6531;
wire n6532;
wire n6533;
wire n6534;
wire n6535;
wire n6536;
wire n6537;
wire n6539;
wire n6540;
wire n6542;
wire n6543;
wire n6544;
wire n6545;
wire n6546;
wire n6547;
wire n6548;
wire n6549;
wire n6550;
wire n6551;
wire n6552;
wire n6553;
wire n6555;
wire n6556;
wire n6557;
wire n6558;
wire n6559;
wire n6560;
wire n6561;
wire n6562;
wire n6563;
wire n6564;
wire n6565;
wire n6566;
wire n6567;
wire n6568;
wire n6569;
wire n6570;
wire n6571;
wire n6572;
wire n6573;
wire n6574;
wire n6577;
wire n6578;
wire n6579;
wire n6580;
wire n6581;
wire n6582;
wire n6583;
wire n6584;
wire n6585;
wire n6587;
wire n6588;
wire n6589;
wire n6590;
wire n6591;
wire n6592;
wire n6593;
wire n6594;
wire n6595;
wire n6599;
wire n6600;
wire n6601;
wire n6602;
wire n6603;
wire n6604;
wire n6605;
wire n6606;
wire n6607;
wire n6608;
wire n6609;
wire n6610;
wire n6611;
wire n6612;
wire n6613;
wire n6614;
wire n6615;
wire n6616;
wire n6617;
wire n6619;
wire n6620;
wire n6621;
wire n6622;
wire n6623;
wire n6624;
wire n6625;
wire n6626;
wire n6627;
wire n6628;
wire n6629;
wire n6630;
wire n6631;
wire n6632;
wire n6633;
wire n6634;
wire n6635;
wire n6636;
wire n6637;
wire n6638;
wire n6639;
wire n6640;
wire n6641;
wire n6642;
wire n6643;
wire n6644;
wire n6646;
wire n6647;
wire n6649;
wire n6650;
wire n6651;
wire n6652;
wire n6653;
wire n6654;
wire n6655;
wire n6656;
wire n6657;
wire n6658;
wire n6659;
wire n6660;
wire n6661;
wire n6662;
wire n6663;
wire n6665;
wire n6666;
wire n6668;
wire n6669;
wire n6670;
wire n6671;
wire n6673;
wire n6674;
wire n6675;
wire n6677;
wire n6678;
wire n6679;
wire n6681;
wire n6682;
wire n6683;
wire n6684;
wire n6685;
wire n6687;
wire n6688;
wire n6689;
wire n6690;
wire n6692;
wire n6693;
wire n6694;
wire n6695;
wire n6696;
wire n6697;
wire n6698;
wire n6701;
wire n6702;
wire n6703;
wire n6704;
wire n6705;
wire n6706;
wire n6707;
wire n6708;
wire n6709;
wire n6710;
wire n6712;
wire n6713;
wire n6714;
wire n6715;
wire n6716;
wire n6717;
wire n6718;
wire n6721;
wire n6722;
wire n6723;
wire n6724;
wire n6725;
wire n6726;
wire n6727;
wire n6728;
wire n6729;
wire n6730;
wire n6731;
wire n6732;
wire n6733;
wire n6734;
wire n6735;
wire n6737;
wire n6738;
wire n6739;
wire n6740;
wire n6741;
wire n6742;
wire n6743;
wire n6744;
wire n6745;
wire n6746;
wire n6747;
wire n6748;
wire n6749;
wire n6750;
wire n6751;
wire n6752;
wire n6753;
wire n6754;
wire n6756;
wire n6757;
wire n6758;
wire n6759;
wire n6760;
wire n6761;
wire n6762;
wire n6763;
wire n6764;
wire n6765;
wire n6766;
wire n6767;
wire n6768;
wire n6769;
wire n6770;
wire n6771;
wire n6773;
wire n6774;
wire n6775;
wire n6776;
wire n6777;
wire n6778;
wire n6779;
wire n6780;
wire n6781;
wire n6782;
wire n6783;
wire n6784;
wire n6785;
wire n6786;
wire n6787;
wire n6788;
wire n6789;
wire n6790;
wire n6792;
wire n6793;
wire n6794;
wire n6795;
wire n6796;
wire n6797;
wire n6798;
wire n6799;
wire n6800;
wire n6801;
wire n6802;
wire n6803;
wire n6804;
wire n6805;
wire n6806;
wire n6807;
wire n6808;
wire n6809;
wire n6810;
wire n6812;
wire n6813;
wire n6815;
wire n6816;
wire n6817;
wire n6818;
wire n6819;
wire n6820;
wire n6821;
wire n6822;
wire n6823;
wire n6826;
wire n6827;
wire n6828;
wire n6829;
wire n6830;
wire n6831;
wire n6832;
wire n6833;
wire n6834;
wire n6835;
wire n6836;
wire n6837;
wire n6838;
wire n6839;
wire n6840;
wire n6841;
wire n6842;
wire n6843;
wire n6844;
wire n6845;
wire n6846;
wire n6847;
wire n6849;
wire n6850;
wire n6851;
wire n6852;
wire n6853;
wire n6854;
wire n6855;
wire n6856;
wire n6858;
wire n6859;
wire n6860;
wire n6861;
wire n6862;
wire n6863;
wire n6864;
wire n6865;
wire n6866;
wire n6867;
wire n6869;
wire n6872;
wire n6873;
wire n6874;
wire n6875;
wire n6876;
wire n6877;
wire n6878;
wire n6879;
wire n6880;
wire n6881;
wire n6882;
wire n6883;
wire n6884;
wire n6885;
wire n6886;
wire n6887;
wire n6888;
wire n6889;
wire n6890;
wire n6891;
wire n6892;
wire n6893;
wire n6894;
wire n6895;
wire n6896;
wire n6897;
wire n6898;
wire n6899;
wire n6900;
wire n6901;
wire n6902;
wire n6903;
wire n6904;
wire n6905;
wire n6906;
wire n6907;
wire n6908;
wire n6909;
wire n6910;
wire n6911;
wire n6912;
wire n6913;
wire n6914;
wire n6915;
wire n6916;
wire n6917;
wire n6918;
wire n6919;
wire n6920;
wire n6921;
wire n6922;
wire n6923;
wire n6924;
wire n6925;
wire n6927;
wire n6928;
wire n6929;
wire n6930;
wire n6931;
wire n6932;
wire n6933;
wire n6934;
wire n6935;
wire n6936;
wire n6937;
wire n6938;
wire n6939;
wire n6940;
wire n6941;
wire n6943;
wire n6944;
wire n6945;
wire n6946;
wire n6947;
wire n6948;
wire n6949;
wire n6951;
wire n6952;
wire n6953;
wire n6954;
wire n6955;
wire n6956;
wire n6957;
wire n6958;
wire n6959;
wire n6960;
wire n6961;
wire n6962;
wire n6963;
wire n6964;
wire n6965;
wire n6966;
wire n6967;
wire n6968;
wire n6969;
wire n6970;
wire n6971;
wire n6972;
wire n6973;
wire n6974;
wire n6975;
wire n6976;
wire n6977;
wire n6978;
wire n6979;
wire n6980;
wire n6981;
wire n6982;
wire n6984;
wire n6985;
wire n6986;
wire n6987;
wire n6988;
wire n6989;
wire n6990;
wire n6992;
wire n6993;
wire n6994;
wire n6995;
wire n6996;
wire n6997;
wire n6998;
wire n6999;
wire n7000;
wire n7001;
wire n7002;
wire n7003;
wire n7004;
wire n7005;
wire n7006;
wire n7007;
wire n7008;
wire n7009;
wire n7010;
wire n7011;
wire n7012;
wire n7014;
wire n7015;
wire n7016;
wire n7017;
wire n7018;
wire n7019;
wire n7020;
wire n7021;
wire n7022;
wire n7023;
wire n7024;
wire n7025;
wire n7026;
wire n7027;
wire n7028;
wire n7029;
wire n7030;
wire n7031;
wire n7032;
wire n7033;
wire n7034;
wire n7035;
wire n7036;
wire n7037;
wire n7038;
wire n7039;
wire n7040;
wire n7041;
wire n7042;
wire n7043;
wire n7044;
wire n7045;
wire n7046;
wire n7047;
wire n7048;
wire n7050;
wire n7051;
wire n7052;
wire n7053;
wire n7055;
wire n7056;
wire n7057;
wire n7058;
wire n7059;
wire n7060;
wire n7062;
wire n7063;
wire n7064;
wire n7065;
wire n7068;
wire n7069;
wire n7070;
wire n7072;
wire n7073;
wire n7074;
wire n7075;
wire n7076;
wire n7077;
wire n7078;
wire n7079;
wire n7080;
wire n7081;
wire n7082;
wire n7083;
wire n7084;
wire n7086;
wire n7087;
wire n7088;
wire n7090;
wire n7091;
wire n7092;
wire n7093;
wire n7094;
wire n7095;
wire n7096;
wire n7097;
wire n7098;
wire n7099;
wire n7100;
wire n7101;
wire n7102;
wire n7103;
wire n7104;
wire n7105;
wire n7108;
wire n7109;
wire n7110;
wire n7111;
wire n7112;
wire n7113;
wire n7114;
wire n7115;
wire n7116;
wire n7118;
wire n7119;
wire n7120;
wire n7121;
wire n7122;
wire n7123;
wire n7124;
wire n7125;
wire n7126;
wire n7127;
wire n7128;
wire n7129;
wire n7131;
wire n7132;
wire n7133;
wire n7134;
wire n7135;
wire n7138;
wire n7139;
wire n7140;
wire n7142;
wire n7143;
wire n7144;
wire n7145;
wire n7146;
wire n7147;
wire n7148;
wire n7149;
wire n7150;
wire n7151;
wire n7152;
wire n7153;
wire n7154;
wire n7155;
wire n7156;
wire n7157;
wire n7158;
wire n7160;
wire n7161;
wire n7162;
wire n7163;
wire n7165;
wire n7166;
wire n7167;
wire n7168;
wire n7169;
wire n7170;
wire n7171;
wire n7172;
wire n7173;
wire n7174;
wire n7175;
wire n7176;
wire n7177;
wire n7178;
wire n7179;
wire n7180;
wire n7181;
wire n7182;
wire n7183;
wire n7184;
wire n7185;
wire n7186;
wire n7187;
wire n7188;
wire n7189;
wire n7190;
wire n7191;
wire n7193;
wire n7194;
wire n7195;
wire n7196;
wire n7197;
wire n7198;
wire n7199;
wire n7200;
wire n7201;
wire n7202;
wire n7203;
wire n7204;
wire n7205;
wire n7206;
wire n7207;
wire n7208;
wire n7209;
wire n7210;
wire n7211;
wire n7212;
wire n7213;
wire n7214;
wire n7215;
wire n7216;
wire n7217;
wire n7218;
wire n7219;
wire n7220;
wire n7221;
wire n7222;
wire n7223;
wire n7224;
wire n7225;
wire n7226;
wire n7228;
wire n7229;
wire n7230;
wire n7231;
wire n7232;
wire n7233;
wire n7234;
wire n7235;
wire n7236;
wire n7237;
wire n7238;
wire n7239;
wire n7240;
wire n7241;
wire n7242;
wire n7243;
wire n7244;
wire n7245;
wire n7246;
wire n7247;
wire n7248;
wire n7249;
wire n7250;
wire n7251;
wire n7252;
wire n7253;
wire n7254;
wire n7255;
wire n7256;
wire n7257;
wire n7258;
wire n7259;
wire n7260;
wire n7261;
wire n7262;
wire n7263;
wire n7264;
wire n7265;
wire n7266;
wire n7267;
wire n7268;
wire n7269;
wire n7270;
wire n7271;
wire n7272;
wire n7273;
wire n7274;
wire n7275;
wire n7276;
wire n7277;
wire n7278;
wire n7279;
wire n7280;
wire n7281;
wire n7282;
wire n7283;
wire n7284;
wire n7286;
wire n7287;
wire n7288;
wire n7289;
wire n7290;
wire n7291;
wire n7292;
wire n7293;
wire n7294;
wire n7295;
wire n7296;
wire n7299;
wire n7300;
wire n7301;
wire n7302;
wire n7303;
wire n7304;
wire n7305;
wire n7306;
wire n7307;
wire n7309;
wire n7310;
wire n7311;
wire n7312;
wire n7313;
wire n7314;
wire n7316;
wire n7317;
wire n7318;
wire n7319;
wire n7320;
wire n7322;
wire n7323;
wire n7324;
wire n7326;
wire n7327;
wire n7328;
wire n7329;
wire n7330;
wire n7331;
wire n7332;
wire n7333;
wire n7334;
wire n7335;
wire n7336;
wire n7337;
wire n7338;
wire n7340;
wire n7341;
wire n7343;
wire n7344;
wire n7345;
wire n7346;
wire n7347;
wire n7348;
wire n7349;
wire n7350;
wire n7351;
wire n7352;
wire n7353;
wire n7354;
wire n7355;
wire n7356;
wire n7357;
wire n7358;
wire n7359;
wire n7360;
wire n7361;
wire n7362;
wire n7363;
wire n7364;
wire n7365;
wire n7366;
wire n7367;
wire n7368;
wire n7369;
wire n7370;
wire n7371;
wire n7372;
wire n7373;
wire n7374;
wire n7375;
wire n7376;
wire n7377;
wire n7378;
wire n7379;
wire n7380;
wire n7381;
wire n7382;
wire n7383;
wire n7384;
wire n7386;
wire n7387;
wire n7388;
wire n7389;
wire n7390;
wire n7391;
wire n7392;
wire n7393;
wire n7394;
wire n7395;
wire n7396;
wire n7397;
wire n7398;
wire n7399;
wire n7400;
wire n7401;
wire n7402;
wire n7403;
wire n7404;
wire n7405;
wire n7406;
wire n7407;
wire n7408;
wire n7409;
wire n7410;
wire n7411;
wire n7412;
wire n7413;
wire n7414;
wire n7415;
wire n7416;
wire n7417;
wire n7418;
wire n7420;
wire n7421;
wire n7423;
wire n7424;
wire n7426;
wire n7427;
wire n7428;
wire n7429;
wire n7431;
wire n7432;
wire n7433;
wire n7434;
wire n7435;
wire n7436;
wire n7437;
wire n7438;
wire n7439;
wire n7440;
wire n7441;
wire n7442;
wire n7443;
wire n7444;
wire n7445;
wire n7446;
wire n7447;
wire n7448;
wire n7449;
wire n7450;
wire n7451;
wire n7452;
wire n7453;
wire n7454;
wire n7455;
wire n7456;
wire n7457;
wire n7458;
wire n7459;
wire n7460;
wire n7461;
wire n7462;
wire n7463;
wire n7464;
wire n7465;
wire n7466;
wire n7467;
wire n7468;
wire n7469;
wire n7470;
wire n7471;
wire n7472;
wire n7473;
wire n7474;
wire n7475;
wire n7476;
wire n7477;
wire n7478;
wire n7479;
wire n7480;
wire n7481;
wire n7482;
wire n7483;
wire n7484;
wire n7485;
wire n7486;
wire n7487;
wire n7488;
wire n7489;
wire n7490;
wire n7491;
wire n7492;
wire n7493;
wire n7494;
wire n7495;
wire n7496;
wire n7497;
wire n7498;
wire n7499;
wire n7500;
wire n7501;
wire n7502;
wire n7504;
wire n7505;
wire n7506;
wire n7507;
wire n7508;
wire n7509;
wire n7510;
wire n7511;
wire n7512;
wire n7513;
wire n7514;
wire n7515;
wire n7516;
wire n7517;
wire n7518;
wire n7519;
wire n7520;
wire n7521;
wire n7522;
wire n7523;
wire n7524;
wire n7525;
wire n7526;
wire n7527;
wire n7528;
wire n7529;
wire n7530;
wire n7531;
wire n7532;
wire n7533;
wire n7534;
wire n7535;
wire n7536;
wire n7537;
wire n7538;
wire n7539;
wire n7540;
wire n7541;
wire n7542;
wire n7543;
wire n7544;
wire n7545;
wire n7546;
wire n7547;
wire n7548;
wire n7549;
wire n7550;
wire n7551;
wire n7552;
wire n7553;
wire n7554;
wire n7555;
wire n7556;
wire n7557;
wire n7558;
wire n7559;
wire n7560;
wire n7561;
wire n7562;
wire n7563;
wire n7564;
wire n7565;
wire n7566;
wire n7567;
wire n7568;
wire n7569;
wire n7570;
wire n7571;
wire n7572;
wire n7573;
wire n7574;
wire n7575;
wire n7576;
wire n7577;
wire n7578;
wire n7579;
wire n7580;
wire n7581;
wire n7582;
wire n7583;
wire n7584;
wire n7585;
wire n7586;
wire n7587;
wire n7588;
wire n7589;
wire n7590;
wire n7591;
wire n7592;
wire n7593;
wire n7594;
wire n7595;
wire n7596;
wire n7597;
wire n7598;
wire n7599;
wire n7600;
wire n7601;
wire n7602;
wire n7603;
wire n7604;
wire n7605;
wire n7606;
wire n7607;
wire n7609;
wire n7610;
wire n7611;
wire n7612;
wire n7613;
wire n7614;
wire n7615;
wire n7616;
wire n7617;
wire n7618;
wire n7619;
wire n7620;
wire n7621;
wire n7622;
wire n7623;
wire n7624;
wire n7625;
wire n7626;
wire n7627;
wire n7628;
wire n7629;
wire n7630;
wire n7631;
wire n7632;
wire n7633;
wire n7634;
wire n7635;
wire n7636;
wire n7637;
wire n7639;
wire n7640;
wire n7641;
wire n7642;
wire n7643;
wire n7644;
wire n7645;
wire n7646;
wire n7648;
wire n7649;
wire n7651;
wire n7653;
wire n7654;
wire n7656;
wire n7657;
wire n7658;
wire n7659;
wire n7660;
wire n7661;
wire n7662;
wire n7663;
wire n7664;
wire n7665;
wire n7666;
wire n7667;
wire n7668;
wire n7669;
wire n7670;
wire n7671;
wire n7673;
wire n7674;
wire n7675;
wire n7677;
wire n7678;
wire n7679;
wire n7680;
wire n7681;
wire n7683;
wire n7684;
wire n7685;
wire n7687;
wire n7688;
wire n7689;
wire n7690;
wire n7691;
wire n7692;
wire n7693;
wire n7694;
wire n7695;
wire n7696;
wire n7697;
wire n7698;
wire n7699;
wire n7700;
wire n7701;
wire n7702;
wire n7703;
wire n7704;
wire n7705;
wire n7706;
wire n7707;
wire n7708;
wire n7709;
wire n7710;
wire n7711;
wire n7712;
wire n7713;
wire n7714;
wire n7715;
wire n7716;
wire n7717;
wire n7718;
wire n7719;
wire n7720;
wire n7721;
wire n7722;
wire n7723;
wire n7724;
wire n7725;
wire n7726;
wire n7727;
wire n7728;
wire n7729;
wire n7730;
wire n7731;
wire n7732;
wire n7733;
wire n7734;
wire n7735;
wire n7736;
wire n7737;
wire n7738;
wire n7739;
wire n7740;
wire n7741;
wire n7743;
wire n7744;
wire n7745;
wire n7746;
wire n7747;
wire n7749;
wire n7750;
wire n7751;
wire n7752;
wire n7753;
wire n7754;
wire n7755;
wire n7756;
wire n7757;
wire n7758;
wire n7760;
wire n7761;
wire n7762;
wire n7763;
wire n7764;
wire n7765;
wire n7766;
wire n7767;
wire n7768;
wire n7770;
wire n7771;
wire n7772;
wire n7773;
wire n7774;
wire n7775;
wire n7776;
wire n7777;
wire n7778;
wire n7779;
wire n7780;
wire n7781;
wire n7782;
wire n7783;
wire n7784;
wire n7785;
wire n7786;
wire n7787;
wire n7788;
wire n7789;
wire n7790;
wire n7791;
wire n7792;
wire n7793;
wire n7794;
wire n7795;
wire n7796;
wire n7798;
wire n7799;
wire n7800;
wire n7802;
wire n7804;
wire n7805;
wire n7807;
wire n7808;
wire n7809;
wire n7810;
wire n7811;
wire n7812;
wire n7813;
wire n7814;
wire n7815;
wire n7816;
wire n7817;
wire n7818;
wire n7820;
wire n7821;
wire n7822;
wire n7823;
wire n7824;
wire n7825;
wire n7826;
wire n7828;
wire n7829;
wire n7830;
wire n7831;
wire n7832;
wire n7833;
wire n7834;
wire n7835;
wire n7836;
wire n7837;
wire n7838;
wire n7841;
wire n7842;
wire n7843;
wire n7844;
wire n7845;
wire n7846;
wire n7847;
wire n7848;
wire n7849;
wire n7850;
wire n7851;
wire n7852;
wire n7854;
wire n7855;
wire n7856;
wire n7857;
wire n7858;
wire n7859;
wire n7860;
wire n7861;
wire n7862;
wire n7863;
wire n7864;
wire n7865;
wire n7866;
wire n7867;
wire n7868;
wire n7870;
wire n7871;
wire n7872;
wire n7873;
wire n7875;
wire n7876;
wire n7877;
wire n7878;
wire n7879;
wire n7880;
wire n7881;
wire n7882;
wire n7883;
wire n7884;
wire n7885;
wire n7886;
wire n7887;
wire n7888;
wire n7889;
wire n7890;
wire n7891;
wire n7892;
wire n7894;
wire n7895;
wire n7896;
wire n7897;
wire n7898;
wire n7899;
wire n7900;
wire n7901;
wire n7902;
wire n7903;
wire n7904;
wire n7905;
wire n7907;
wire n7908;
wire n7909;
wire n7910;
wire n7912;
wire n7913;
wire n7914;
wire n7915;
wire n7916;
wire n7917;
wire n7918;
wire n7919;
wire n7920;
wire n7921;
wire n7922;
wire n7923;
wire n7924;
wire n7925;
wire n7926;
wire n7927;
wire n7928;
wire n7929;
wire n7930;
wire n7931;
wire n7932;
wire n7933;
wire n7934;
wire n7935;
wire n7936;
wire n7938;
wire n7939;
wire n7940;
wire n7941;
wire n7942;
wire n7943;
wire n7944;
wire n7945;
wire n7946;
wire n7947;
wire n7948;
wire n7949;
wire n7950;
wire n7951;
wire n7952;
wire n7953;
wire n7954;
wire n7955;
wire n7956;
wire n7957;
wire n7958;
wire n7959;
wire n7960;
wire n7961;
wire n7962;
wire n7963;
wire n7964;
wire n7965;
wire n7966;
wire n7967;
wire n7968;
wire n7969;
wire n7970;
wire n7971;
wire n7972;
wire n7973;
wire n7974;
wire n7975;
wire n7976;
wire n7977;
wire n7978;
wire n7979;
wire n7980;
wire n7981;
wire n7982;
wire n7983;
wire n7985;
wire n7986;
wire n7987;
wire n7988;
wire n7989;
wire n7990;
wire n7991;
wire n7992;
wire n7993;
wire n7994;
wire n7995;
wire n7996;
wire n7997;
wire n7998;
wire n7999;
wire n8000;
wire n8001;
wire n8002;
wire n8003;
wire n8004;
wire n8005;
wire n8006;
wire n8007;
wire n8008;
wire n8009;
wire n8010;
wire n8011;
wire n8012;
wire n8013;
wire n8014;
wire n8015;
wire n8016;
wire n8017;
wire n8018;
wire n8019;
wire n8020;
wire n8021;
wire n8022;
wire n8023;
wire n8024;
wire n8025;
wire n8026;
wire n8027;
wire n8028;
wire n8029;
wire n8030;
wire n8031;
wire n8032;
wire n8033;
wire n8034;
wire n8035;
wire n8036;
wire n8037;
wire n8038;
wire n8039;
wire n8040;
wire n8041;
wire n8042;
wire n8043;
wire n8044;
wire n8045;
wire n8047;
wire n8048;
wire n8049;
wire n8050;
wire n8051;
wire n8052;
wire n8053;
wire n8054;
wire n8055;
wire n8056;
wire n8057;
wire n8058;
wire n8059;
wire n8060;
wire n8061;
wire n8062;
wire n8063;
wire n8064;
wire n8067;
wire n8068;
wire n8069;
wire n8072;
wire n8073;
wire n8074;
wire n8075;
wire n8076;
wire n8077;
wire n8078;
wire n8079;
wire n8080;
wire n8081;
wire n8082;
wire n8083;
wire n8084;
wire n8085;
wire n8086;
wire n8087;
wire n8088;
wire n8089;
wire n8090;
wire n8091;
wire n8092;
wire n8093;
wire n8094;
wire n8095;
wire n8096;
wire n8097;
wire n8098;
wire n8099;
wire n8100;
wire n8101;
wire n8102;
wire n8103;
wire n8104;
wire n8105;
wire n8106;
wire n8107;
wire n8108;
wire n8109;
wire n8110;
wire n8111;
wire n8113;
wire n8114;
wire n8115;
wire n8116;
wire n8117;
wire n8118;
wire n8119;
wire n8120;
wire n8121;
wire n8122;
wire n8123;
wire n8124;
wire n8125;
wire n8126;
wire n8127;
wire n8128;
wire n8129;
wire n8130;
wire n8131;
wire n8132;
wire n8133;
wire n8134;
wire n8135;
wire n8136;
wire n8137;
wire n8138;
wire n8139;
wire n8140;
wire n8141;
wire n8142;
wire n8143;
wire n8144;
wire n8145;
wire n8146;
wire n8147;
wire n8148;
wire n8149;
wire n8150;
wire n8151;
wire n8152;
wire n8153;
wire n8154;
wire n8155;
wire n8156;
wire n8157;
wire n8158;
wire n8159;
wire n8160;
wire n8161;
wire n8162;
wire n8163;
wire n8164;
wire n8165;
wire n8166;
wire n8167;
wire n8168;
wire n8169;
wire n8170;
wire n8171;
wire n8172;
wire n8173;
wire n8174;
wire n8175;
wire n8176;
wire n8177;
wire n8178;
wire n8179;
wire n8180;
wire n8181;
wire n8182;
wire n8183;
wire n8184;
wire n8185;
wire n8186;
wire n8187;
wire n8188;
wire n8189;
wire n8190;
wire n8191;
wire n8192;
wire n8193;
wire n8194;
wire n8195;
wire n8196;
wire n8197;
wire n8198;
wire n8199;
wire n8200;
wire n8201;
wire n8202;
wire n8203;
wire n8204;
wire n8205;
wire n8206;
wire n8207;
wire n8208;
wire n8209;
wire n8210;
wire n8211;
wire n8212;
wire n8213;
wire n8214;
wire n8215;
wire n8216;
wire n8217;
wire n8218;
wire n8219;
wire n8220;
wire n8221;
wire n8222;
wire n8223;
wire n8224;
wire n8225;
wire n8226;
wire n8227;
wire n8228;
wire n8229;
wire n8230;
wire n8231;
wire n8232;
wire n8233;
wire n8234;
wire n8235;
wire n8236;
wire n8237;
wire n8238;
wire n8239;
wire n8240;
wire n8241;
wire n8242;
wire n8243;
wire n8244;
wire n8245;
wire n8246;
wire n8247;
wire n8248;
wire n8249;
wire n8250;
wire n8251;
wire n8252;
wire n8253;
wire n8254;
wire n8255;
wire n8256;
wire n8257;
wire n8258;
wire n8259;
wire n8260;
wire n8261;
wire n8262;
wire n8263;
wire n8264;
wire n8265;
wire n8266;
wire n8267;
wire n8268;
wire n8269;
wire n8270;
wire n8271;
wire n8272;
wire n8273;
wire n8274;
wire n8275;
wire n8276;
wire n8277;
wire n8278;
wire n8279;
wire n8280;
wire n8281;
wire n8282;
wire n8283;
wire n8284;
wire n8285;
wire n8286;
wire n8287;
wire n8288;
wire n8289;
wire n8290;
wire n8291;
wire n8292;
wire n8293;
wire n8294;
wire n8295;
wire n8296;
wire n8297;
wire n8298;
wire n8299;
wire n8300;
wire n8301;
wire n8302;
wire n8303;
wire n8304;
wire n8305;
wire n8306;
wire n8307;
wire n8308;
wire n8309;
wire n8310;
wire n8311;
wire n8312;
wire n8313;
wire n8315;
wire n8316;
wire n8317;
wire n8318;
wire n8319;
wire n8320;
wire n8321;
wire n8322;
wire n8323;
wire n8324;
wire n8325;
wire n8326;
wire n8327;
wire n8328;
wire n8329;
wire n8330;
wire n8331;
wire n8332;
wire n8333;
wire n8334;
wire n8335;
wire n8336;
wire n8337;
wire n8338;
wire n8339;
wire n8340;
wire n8341;
wire n8342;
wire n8343;
wire n8344;
wire n8345;
wire n8346;
wire n8347;
wire n8348;
wire n8350;
wire n8351;
wire n8352;
wire n8353;
wire n8354;
wire n8355;
wire n8356;
wire n8357;
wire n8358;
wire n8359;
wire n8360;
wire n8361;
wire n8362;
wire n8363;
wire n8364;
wire n8365;
wire n8366;
wire n8367;
wire n8369;
wire n8370;
wire n8371;
wire n8372;
wire n8373;
wire n8374;
wire n8375;
wire n8376;
wire n8377;
wire n8378;
wire n8379;
wire n8380;
wire n8381;
wire n8382;
wire n8383;
wire n8384;
wire n8385;
wire n8386;
wire n8387;
wire n8388;
wire n8389;
wire n8390;
wire n8391;
wire n8392;
wire n8393;
wire n8394;
wire n8395;
wire n8396;
wire n8397;
wire n8398;
wire n8399;
wire n8400;
wire n8401;
wire n8402;
wire n8403;
wire n8404;
wire n8405;
wire n8406;
wire n8407;
wire n8408;
wire n8409;
wire n8410;
wire n8411;
wire n8412;
wire n8413;
wire n8414;
wire n8415;
wire n8416;
wire n8417;
wire n8418;
wire n8419;
wire n8420;
wire n8421;
wire n8422;
wire n8423;
wire n8424;
wire n8425;
wire n8426;
wire n8427;
wire n8428;
wire n8429;
wire n8430;
wire n8431;
wire n8432;
wire n8433;
wire n8434;
wire n8435;
wire n8436;
wire n8437;
wire n8438;
wire n8439;
wire n8440;
wire n8442;
wire n8443;
wire n8444;
wire n8445;
wire n8446;
wire n8447;
wire n8448;
wire n8449;
wire n8450;
wire n8451;
wire n8452;
wire n8453;
wire n8454;
wire n8455;
wire n8456;
wire n8457;
wire n8458;
wire n8459;
wire n8460;
wire n8461;
wire n8462;
wire n8463;
wire n8465;
wire n8466;
wire n8467;
wire n8468;
wire n8469;
wire n8470;
wire n8471;
wire n8472;
wire n8473;
wire n8474;
wire n8475;
wire n8476;
wire n8477;
wire n8478;
wire n8479;
wire n8480;
wire n8481;
wire n8482;
wire n8483;
wire n8484;
wire n8486;
wire n8487;
wire n8488;
wire n8489;
wire n8490;
wire n8491;
wire n8492;
wire n8493;
wire n8494;
wire n8495;
wire n8496;
wire n8497;
wire n8498;
wire n8499;
wire n8500;
wire n8501;
wire n8502;
wire n8503;
wire n8504;
wire n8505;
wire n8506;
wire n8507;
wire n8508;
wire n8509;
wire n8510;
wire n8511;
wire n8512;
wire n8513;
wire n8514;
wire n8515;
wire n8516;
wire n8517;
wire n8518;
wire n8519;
wire n8520;
wire n8521;
wire n8522;
wire n8523;
wire n8524;
wire n8525;
wire n8526;
wire n8527;
wire n8528;
wire n8529;
wire n8530;
wire n8531;
wire n8532;
wire n8533;
wire n8534;
wire n8535;
wire n8537;
wire n8538;
wire n8539;
wire n8540;
wire n8541;
wire n8542;
wire n8543;
wire n8544;
wire n8545;
wire n8546;
wire n8547;
wire n8548;
wire n8549;
wire n8550;
wire n8551;
wire n8553;
wire n8554;
wire n8555;
wire n8556;
wire n8557;
wire n8558;
wire n8559;
wire n8560;
wire n8561;
wire n8562;
wire n8563;
wire n8564;
wire n8565;
wire n8566;
wire n8567;
wire n8568;
wire n8569;
wire n8570;
wire n8571;
wire n8572;
wire n8573;
wire n8574;
wire n8575;
wire n8576;
wire n8577;
wire n8578;
wire n8579;
wire n8580;
wire n8581;
wire n8582;
wire n8583;
wire n8586;
wire n8587;
wire n8588;
wire n8589;
wire n8590;
wire n8591;
wire n8592;
wire n8593;
wire n8594;
wire n8595;
wire n8596;
wire n8597;
wire n8598;
wire n8599;
wire n8600;
wire n8601;
wire n8602;
wire n8603;
wire n8604;
wire n8605;
wire n8606;
wire n8607;
wire n8608;
wire n8609;
wire n8610;
wire n8611;
wire n8613;
wire n8614;
wire n8615;
wire n8616;
wire n8617;
wire n8618;
wire n8619;
wire n8620;
wire n8621;
wire n8622;
wire n8623;
wire n8624;
wire n8625;
wire n8626;
wire n8627;
wire n8628;
wire n8629;
wire n8630;
wire n8631;
wire n8632;
wire n8633;
wire n8634;
wire n8635;
wire n8636;
wire n8637;
wire n8638;
wire n8639;
wire n8640;
wire n8642;
wire n8643;
wire n8644;
wire n8645;
wire n8646;
wire n8647;
wire n8648;
wire n8649;
wire n8650;
wire n8651;
wire n8652;
wire n8653;
wire n8654;
wire n8655;
wire n8656;
wire n8657;
wire n8658;
wire n8659;
wire n8660;
wire n8661;
wire n8662;
wire n8663;
wire n8664;
wire n8665;
wire n8666;
wire n8667;
wire n8668;
wire n8669;
wire n8670;
wire n8671;
wire n8672;
wire n8673;
wire n8674;
wire n8675;
wire n8676;
wire n8677;
wire n8678;
wire n8679;
wire n8680;
wire n8681;
wire n8682;
wire n8683;
wire n8684;
wire n8685;
wire n8686;
wire n8687;
wire n8688;
wire n8689;
wire n8690;
wire n8691;
wire n8692;
wire n8693;
wire n8694;
wire n8695;
wire n8696;
wire n8697;
wire n8698;
wire n8699;
wire n8700;
wire n8701;
wire n8702;
wire n8703;
wire n8704;
wire n8705;
wire n8706;
wire n8707;
wire n8708;
wire n8709;
wire n8710;
wire n8711;
wire n8712;
wire n8713;
wire n8714;
wire n8715;
wire n8716;
wire n8717;
wire n8718;
wire n8719;
wire n8720;
wire n8721;
wire n8722;
wire n8723;
wire n8724;
wire n8725;
wire n8726;
wire n8727;
wire n8728;
wire n8729;
wire n8730;
wire n8731;
wire n8732;
wire n8733;
wire n8734;
wire n8735;
wire n8736;
wire n8737;
wire n8738;
wire n8739;
wire n8740;
wire n8741;
wire n8742;
wire n8743;
wire n8745;
wire n8746;
wire n8747;
wire n8748;
wire n8749;
wire n8750;
wire n8751;
wire n8752;
wire n8753;
wire n8754;
wire n8755;
wire n8756;
wire n8757;
wire n8758;
wire n8759;
wire n8760;
wire n8761;
wire n8762;
wire n8763;
wire n8764;
wire n8765;
wire n8766;
wire n8767;
wire n8768;
wire n8769;
wire n8770;
wire n8771;
wire n8772;
wire n8773;
wire n8774;
wire n8775;
wire n8776;
wire n8777;
wire n8778;
wire n8779;
wire n8780;
wire n8781;
wire n8782;
wire n8783;
wire n8784;
wire n8785;
wire n8786;
wire n8787;
wire n8788;
wire n8789;
wire n8790;
wire n8791;
wire n8792;
wire n8793;
wire n8794;
wire n8795;
wire n8796;
wire n8797;
wire n8798;
wire n8799;
wire n8800;
wire n8801;
wire n8802;
wire n8803;
wire n8804;
wire n8805;
wire n8806;
wire n8807;
wire n8808;
wire n8809;
wire n8810;
wire n8811;
wire n8812;
wire n8813;
wire n8814;
wire n8815;
wire n8816;
wire n8817;
wire n8818;
wire n8819;
wire n8820;
wire n8821;
wire n8822;
wire n8823;
wire n8824;
wire n8825;
wire n8826;
wire n8827;
wire n8828;
wire n8829;
wire n8830;
wire n8831;
wire n8832;
wire n8833;
wire n8834;
wire n8835;
wire n8836;
wire n8837;
wire n8838;
wire n8839;
wire n8840;
wire n8841;
wire n8842;
wire n8843;
wire n8844;
wire n8845;
wire n8846;
wire n8847;
wire n8848;
wire n8849;
wire n8850;
wire n8851;
wire n8852;
wire n8853;
wire n8854;
wire n8855;
wire n8856;
wire n8857;
wire n8858;
wire n8859;
wire n8860;
wire n8862;
wire n8863;
wire n8864;
wire n8865;
wire n8866;
wire n8868;
wire n8869;
wire n8870;
wire n8871;
wire n8872;
wire n8873;
wire n8874;
wire n8875;
wire n8876;
wire n8877;
wire n8878;
wire n8879;
wire n8880;
wire n8881;
wire n8882;
wire n8883;
wire n8884;
wire n8885;
wire n8886;
wire n8887;
wire n8888;
wire n8889;
wire n8890;
wire n8891;
wire n8892;
wire n8893;
wire n8894;
wire n8895;
wire n8896;
wire n8897;
wire n8898;
wire n8899;
wire n8900;
wire n8901;
wire n8902;
wire n8903;
wire n8904;
wire n8906;
wire n8907;
wire n8908;
wire n8909;
wire n8910;
wire n8911;
wire n8912;
wire n8913;
wire n8914;
wire n8915;
wire n8916;
wire n8917;
wire n8918;
wire n8919;
wire n8920;
wire n8921;
wire n8922;
wire n8923;
wire n8924;
wire n8925;
wire n8926;
wire n8927;
wire n8928;
wire n8929;
wire n8930;
wire n8931;
wire n8932;
wire n8933;
wire n8934;
wire n8935;
wire n8936;
wire n8937;
wire n8938;
wire n8939;
wire n8940;
wire n8941;
wire n8942;
wire n8943;
wire n8944;
wire n8945;
wire n8946;
wire n8947;
wire n8948;
wire n8949;
wire n8950;
wire n8951;
wire n8952;
wire n8953;
wire n8954;
wire n8955;
wire n8956;
wire n8957;
wire n8958;
wire n8959;
wire n8960;
wire n8961;
wire n8962;
wire n8963;
wire n8964;
wire n8965;
wire n8966;
wire n8967;
wire n8968;
wire n8969;
wire n8970;
wire n8971;
wire n8972;
wire n8973;
wire n8974;
wire n8975;
wire n8976;
wire n8977;
wire n8978;
wire n8979;
wire n8980;
wire n8981;
wire n8982;
wire n8983;
wire n8984;
wire n8985;
wire n8986;
wire n8987;
wire n8988;
wire n8989;
wire n8990;
wire n8991;
wire n8992;
wire n8993;
wire n8994;
wire n8995;
wire n8996;
wire n8997;
wire n8998;
wire n8999;
wire n9000;
wire n9001;
wire n9003;
wire n9004;
wire n9005;
wire n9006;
wire n9007;
wire n9008;
wire n9009;
wire n9010;
wire n9011;
wire n9012;
wire n9013;
wire n9014;
wire n9015;
wire n9017;
wire n9018;
wire n9019;
wire n9020;
wire n9021;
wire n9022;
wire n9023;
wire n9024;
wire n9025;
wire n9026;
wire n9027;
wire n9028;
wire n9029;
wire n9030;
wire n9031;
wire n9032;
wire n9033;
wire n9034;
wire n9035;
wire n9036;
wire n9037;
wire n9038;
wire n9039;
wire n9040;
wire n9041;
wire n9042;
wire n9043;
wire n9044;
wire n9045;
wire n9046;
wire n9047;
wire n9048;
wire n9049;
wire n9050;
wire n9051;
wire n9052;
wire n9053;
wire n9054;
wire n9055;
wire n9057;
wire n9058;
wire n9059;
wire n9060;
wire n9061;
wire n9062;
wire n9063;
wire n9064;
wire n9065;
wire n9066;
wire n9067;
wire n9068;
wire n9069;
wire n9070;
wire n9071;
wire n9072;
wire n9073;
wire n9074;
wire n9075;
wire n9076;
wire n9077;
wire n9078;
wire n9079;
wire n9080;
wire n9081;
wire n9082;
wire n9084;
wire n9085;
wire n9086;
wire n9087;
wire n9088;
wire n9089;
wire n9090;
wire n9091;
wire n9092;
wire n9093;
wire n9094;
wire n9095;
wire n9096;
wire n9097;
wire n9098;
wire n9099;
wire n9100;
wire n9102;
wire n9103;
wire n9104;
wire n9105;
wire n9106;
wire n9107;
wire n9108;
wire n9109;
wire n9110;
wire n9111;
wire n9112;
wire n9113;
wire n9115;
wire n9116;
wire n9117;
wire n9118;
wire n9119;
wire n9120;
wire n9121;
wire n9122;
wire n9123;
wire n9124;
wire n9125;
wire n9126;
wire n9127;
wire n9128;
wire n9129;
wire n9130;
wire n9131;
wire n9132;
wire n9133;
wire n9135;
wire n9136;
wire n9137;
wire n9138;
wire n9139;
wire n9140;
wire n9141;
wire n9142;
wire n9143;
wire n9144;
wire n9145;
wire n9146;
wire n9147;
wire n9148;
wire n9149;
wire n9150;
wire n9151;
wire n9152;
wire n9153;
wire n9154;
wire n9155;
wire n9156;
wire n9158;
wire n9159;
wire n9160;
wire n9161;
wire n9162;
wire n9163;
wire n9164;
wire n9165;
wire n9166;
wire n9167;
wire n9168;
wire n9169;
wire n9170;
wire n9171;
wire n9172;
wire n9173;
wire n9174;
wire n9175;
wire n9176;
wire n9177;
wire n9178;
wire n9179;
wire n9180;
wire n9181;
wire n9182;
wire n9183;
wire n9184;
wire n9185;
wire n9186;
wire n9187;
wire n9188;
wire n9189;
wire n9190;
wire n9191;
wire n9192;
wire n9193;
wire n9194;
wire n9195;
wire n9196;
wire n9197;
wire n9198;
wire n9199;
wire n9200;
wire n9201;
wire n9202;
wire n9203;
wire n9204;
wire n9205;
wire n9206;
wire n9207;
wire n9208;
wire n9209;
wire n9210;
wire n9211;
wire n9212;
wire n9213;
wire n9214;
wire n9215;
wire n9216;
wire n9217;
wire n9218;
wire n9219;
wire n9220;
wire n9221;
wire n9222;
wire n9223;
wire n9224;
wire n9225;
wire n9226;
wire n9227;
wire n9228;
wire n9229;
wire n9230;
wire n9231;
wire n9232;
wire n9233;
wire n9234;
wire n9235;
wire n9236;
wire n9237;
wire n9238;
wire n9239;
wire n9240;
wire n9241;
wire n9242;
wire n9243;
wire n9245;
wire n9246;
wire n9247;
wire n9248;
wire n9249;
wire n9250;
wire n9251;
wire n9252;
wire n9253;
wire n9254;
wire n9255;
wire n9256;
wire n9257;
wire n9258;
wire n9259;
wire n9260;
wire n9261;
wire n9262;
wire n9263;
wire n9264;
wire n9265;
wire n9266;
wire n9267;
wire n9268;
wire n9269;
wire n9270;
wire n9271;
wire n9272;
wire n9273;
wire n9274;
wire n9275;
wire n9276;
wire n9277;
wire n9278;
wire n9279;
wire n9280;
wire n9281;
wire n9282;
wire n9283;
wire n9284;
wire n9285;
wire n9286;
wire n9287;
wire n9288;
wire n9289;
wire n9290;
wire n9291;
wire n9292;
wire n9293;
wire n9294;
wire n9295;
wire n9296;
wire n9297;
wire n9298;
wire n9299;
wire n9300;
wire n9301;
wire n9302;
wire n9303;
wire n9304;
wire n9305;
wire n9306;
wire n9307;
wire n9308;
wire n9309;
wire n9310;
wire n9311;
wire n9312;
wire n9314;
wire n9315;
wire n9316;
wire n9317;
wire n9318;
wire n9319;
wire n9320;
wire n9321;
wire n9322;
wire n9323;
wire n9324;
wire n9325;
wire n9326;
wire n9327;
wire n9328;
wire n9329;
wire n9330;
wire n9331;
wire n9332;
wire n9333;
wire n9334;
wire n9335;
wire n9336;
wire n9337;
wire n9338;
wire n9339;
wire n9340;
wire n9341;
wire n9342;
wire n9343;
wire n9344;
wire n9345;
wire n9346;
wire n9347;
wire n9348;
wire n9349;
wire n9350;
wire n9351;
wire n9352;
wire n9353;
wire n9354;
wire n9355;
wire n9356;
wire n9357;
wire n9358;
wire n9359;
wire n9360;
wire n9361;
wire n9362;
wire n9363;
wire n9364;
wire n9365;
wire n9366;
wire n9367;
wire n9368;
wire n9369;
wire n9370;
wire n9371;
wire n9372;
wire n9374;
wire n9375;
wire n9376;
wire n9377;
wire n9378;
wire n9379;
wire n9380;
wire n9381;
wire n9382;
wire n9383;
wire n9384;
wire n9385;
wire n9386;
wire n9387;
wire n9388;
wire n9389;
wire n9390;
wire n9391;
wire n9392;
wire n9393;
wire n9394;
wire n9395;
wire n9396;
wire n9397;
wire n9398;
wire n9399;
wire n9400;
wire n9401;
wire n9402;
wire n9403;
wire n9404;
wire n9405;
wire n9406;
wire n9407;
wire n9408;
wire n9409;
wire n9410;
wire n9411;
wire n9412;
wire n9413;
wire n9414;
wire n9415;
wire n9416;
wire n9417;
wire n9418;
wire n9419;
wire n9420;
wire n9421;
wire n9422;
wire n9423;
wire n9424;
wire n9425;
wire n9426;
wire n9427;
wire n9428;
wire n9429;
wire n9430;
wire n9431;
wire n9432;
wire n9433;
wire n9434;
wire n9435;
wire n9436;
wire n9437;
wire n9438;
wire n9439;
wire n9440;
wire n9441;
wire n9442;
wire n9443;
wire n9444;
wire n9445;
wire n9446;
wire n9447;
wire n9448;
wire n9449;
wire n9450;
wire n9451;
wire n9454;
wire n9455;
wire n9456;
wire n9457;
wire n9458;
wire n9459;
wire n9460;
wire n9461;
wire n9462;
wire n9463;
wire n9464;
wire n9465;
wire n9466;
wire n9467;
wire n9468;
wire n9469;
wire n9470;
wire n9471;
wire n9472;
wire n9473;
wire n9474;
wire n9475;
wire n9476;
wire n9477;
wire n9478;
wire n9479;
wire n9480;
wire n9481;
wire n9482;
wire n9483;
wire n9484;
wire n9485;
wire n9486;
wire n9487;
wire n9488;
wire n9489;
wire n9490;
wire n9491;
wire n9492;
wire n9493;
wire n9494;
wire n9495;
wire n9496;
wire n9497;
wire n9498;
wire n9499;
wire n9500;
wire n9501;
wire n9502;
wire n9503;
wire n9504;
wire n9505;
wire n9506;
wire n9507;
wire n9508;
wire n9509;
wire n9510;
wire n9511;
wire n9512;
wire n9513;
wire n9514;
wire n9515;
wire n9516;
wire n9517;
wire n9518;
wire n9519;
wire n9520;
wire n9521;
wire n9522;
wire n9523;
wire n9524;
wire n9525;
wire n9526;
wire n9527;
wire n9528;
wire n9529;
wire n9530;
wire n9531;
wire n9532;
wire n9533;
wire n9534;
wire n9535;
wire n9536;
wire n9537;
wire n9538;
wire n9539;
wire n9540;
wire n9541;
wire n9542;
wire n9543;
wire n9544;
wire n9545;
wire n9546;
wire n9547;
wire n9548;
wire n9549;
wire n9550;
wire n9551;
wire n9552;
wire n9553;
wire n9554;
wire n9555;
wire n9556;
wire n9557;
wire n9558;
wire n9559;
wire n9560;
wire n9561;
wire n9562;
wire n9563;
wire n9564;
wire n9565;
wire n9566;
wire n9567;
wire n9568;
wire n9569;
wire n9570;
wire n9571;
wire n9572;
wire n9573;
wire n9574;
wire n9575;
wire n9576;
wire n9577;
wire n9578;
wire n9579;
wire n9580;
wire n9581;
wire n9582;
wire n9583;
wire n9584;
wire n9585;
wire n9586;
wire n9587;
wire n9588;
wire n9589;
wire n9590;
wire n9591;
wire n9592;
wire n9593;
wire n9594;
wire n9595;
wire n9596;
wire n9597;
wire n9598;
wire n9599;
wire n9600;
wire n9601;
wire n9602;
wire n9603;
wire n9604;
wire n9605;
wire n9606;
wire n9607;
wire n9608;
wire n9609;
wire n9610;
wire n9611;
wire n9612;
wire n9613;
wire n9614;
wire n9615;
wire n9616;
wire n9617;
wire n9618;
wire n9619;
wire n9620;
wire n9621;
wire n9622;
wire n9623;
wire n9624;
wire n9625;
wire n9626;
wire n9627;
wire n9628;
wire n9629;
wire n9630;
wire n9631;
wire n9632;
wire n9635;
wire n9637;
wire n9638;
wire n9639;
wire n9640;
wire n9641;
wire n9642;
wire n9643;
wire n9644;
wire n9645;
wire n9646;
wire n9647;
wire n9648;
wire n9649;
wire n9650;
wire n9651;
wire n9652;
wire n9653;
wire n9654;
wire n9655;
wire n9656;
wire n9657;
wire n9659;
wire n9660;
wire n9661;
wire n9662;
wire n9663;
wire n9664;
wire n9665;
wire n9666;
wire n9667;
wire n9668;
wire n9669;
wire n9670;
wire n9671;
wire n9672;
wire n9673;
wire n9674;
wire n9675;
wire n9676;
wire n9677;
wire n9678;
wire n9679;
wire n9680;
wire n9681;
wire n9682;
wire n9683;
wire n9684;
wire n9685;
wire n9686;
wire n9687;
wire n9688;
wire n9689;
wire n9690;
wire n9691;
wire n9692;
wire n9693;
wire n9694;
wire n9695;
wire n9696;
wire n9697;
wire n9698;
wire n9699;
wire n9700;
wire n9701;
wire n9702;
wire n9703;
wire n9704;
wire n9705;
wire n9706;
wire n9707;
wire n9708;
wire n9709;
wire n9710;
wire n9711;
wire n9713;
wire n9714;
wire n9715;
wire n9716;
wire n9717;
wire n9718;
wire n9719;
wire n9720;
wire n9721;
wire n9722;
wire n9723;
wire n9724;
wire n9725;
wire n9726;
wire n9727;
wire n9728;
wire n9729;
wire n9730;
wire n9731;
wire n9732;
wire n9733;
wire n9735;
wire n9736;
wire n9737;
wire n9738;
wire n9740;
wire n9741;
wire n9742;
wire n9743;
wire n9744;
wire n9745;
wire n9746;
wire n9747;
wire n9748;
wire n9749;
wire n9750;
wire n9751;
wire n9752;
wire n9753;
wire n9754;
wire n9755;
wire n9756;
wire n9757;
wire n9758;
wire n9759;
wire n9760;
wire n9761;
wire n9762;
wire n9765;
wire n9766;
wire n9767;
wire n9768;
wire n9769;
wire n9770;
wire n9771;
wire n9772;
wire n9773;
wire n9774;
wire n9775;
wire n9776;
wire n9777;
wire n9778;
wire n9779;
wire n9780;
wire n9781;
wire n9782;
wire n9783;
wire n9784;
wire n9785;
wire n9786;
wire n9787;
wire n9788;
wire n9789;
wire n9790;
wire n9791;
wire n9792;
wire n9793;
wire n9794;
wire n9795;
wire n9796;
wire n9797;
wire n9798;
wire n9799;
wire n9800;
wire n9801;
wire n9802;
wire n9803;
wire n9804;
wire n9805;
wire n9806;
wire n9807;
wire n9808;
wire n9809;
wire n9810;
wire n9811;
wire n9812;
wire n9813;
wire n9814;
wire n9815;
wire n9816;
wire n9817;
wire n9818;
wire n9819;
wire n9820;
wire n9821;
wire n9822;
wire n9823;
wire n9824;
wire n9825;
wire n9826;
wire n9827;
wire n9828;
wire n9829;
wire n9830;
wire n9831;
wire n9832;
wire n9833;
wire n9834;
wire n9835;
wire n9836;
wire n9837;
wire n9838;
wire n9839;
wire n9840;
wire n9841;
wire n9842;
wire n9843;
wire n9844;
wire n9845;
wire n9846;
wire n9847;
wire n9848;
wire n9849;
wire n9850;
wire n9851;
wire n9852;
wire n9853;
wire n9854;
wire n9855;
wire n9856;
wire n9857;
wire n9858;
wire n9859;
wire n9860;
wire n9861;
wire n9862;
wire n9863;
wire n9864;
wire n9865;
wire n9866;
wire n9867;
wire n9868;
wire n9870;
wire n9871;
wire n9872;
wire n9873;
wire n9874;
wire n9875;
wire n9876;
wire n9877;
wire n9878;
wire n9879;
wire n9880;
wire n9881;
wire n9882;
wire n9883;
wire n9884;
wire n9885;
wire n9886;
wire n9887;
wire n9888;
wire n9889;
wire n9890;
wire n9891;
wire n9892;
wire n9893;
wire n9894;
wire n9895;
wire n9896;
wire n9897;
wire n9898;
wire n9899;
wire n9900;
wire n9901;
wire n9902;
wire n9903;
wire n9904;
wire n9905;
wire n9906;
wire n9907;
wire n9908;
wire n9909;
wire n9910;
wire n9911;
wire n9912;
wire n9913;
wire n9914;
wire n9915;
wire n9916;
wire n9917;
wire n9918;
wire n9919;
wire n9920;
wire n9921;
wire n9923;
wire n9924;
wire n9925;
wire n9926;
wire n9927;
wire n9928;
wire n9929;
wire n9930;
wire n9931;
wire n9932;
wire n9933;
wire n9934;
wire n9935;
wire n9936;
wire n9937;
wire n9938;
wire n9939;
wire n9940;
wire n9941;
wire n9942;
wire n9943;
wire n9944;
wire n9945;
wire n9946;
wire n9947;
wire n9948;
wire n9949;
wire n9950;
wire n9951;
wire n9952;
wire n9953;
wire n9954;
wire n9955;
wire n9956;
wire n9957;
wire n9958;
wire n9959;
wire n9960;
wire n9961;
wire n9962;
wire n9963;
wire n9964;
wire n9965;
wire n9966;
wire n9967;
wire n9968;
wire n9969;
wire n9970;
wire n9971;
wire n9973;
wire n9974;
wire n9975;
wire n9976;
wire n9977;
wire n9978;
wire n9979;
wire n9980;
wire n9981;
wire n9982;
wire n9983;
wire n9984;
wire n9985;
wire n9986;
wire n9987;
wire n9988;
wire n9989;
wire n9990;
wire n9991;
wire n9992;
wire n9993;
wire n9994;
wire n9995;
wire n9996;
wire n9997;
wire n9998;
wire n9999;
wire n10000;
wire n10001;
wire n10002;
wire n10003;
wire n10004;
wire n10005;
wire n10006;
wire n10007;
wire n10008;
wire n10009;
wire n10010;
wire n10011;
wire n10012;
wire n10013;
wire n10014;
wire n10015;
wire n10016;
wire n10017;
wire n10018;
wire n10019;
wire n10020;
wire n10021;
wire n10022;
wire n10023;
wire n10024;
wire n10025;
wire n10026;
wire n10027;
wire n10028;
wire n10029;
wire n10030;
wire n10031;
wire n10032;
wire n10033;
wire n10034;
wire n10035;
wire n10036;
wire n10037;
wire n10038;
wire n10040;
wire n10041;
wire n10042;
wire n10043;
wire n10044;
wire n10045;
wire n10046;
wire n10047;
wire n10048;
wire n10049;
wire n10050;
wire n10051;
wire n10052;
wire n10053;
wire n10054;
wire n10055;
wire n10056;
wire n10057;
wire n10058;
wire n10059;
wire n10060;
wire n10061;
wire n10062;
wire n10063;
wire n10064;
wire n10065;
wire n10066;
wire n10067;
wire n10068;
wire n10069;
wire n10070;
wire n10071;
wire n10073;
wire n10074;
wire n10075;
wire n10076;
wire n10077;
wire n10078;
wire n10079;
wire n10080;
wire n10081;
wire n10082;
wire n10083;
wire n10084;
wire n10085;
wire n10086;
wire n10087;
wire n10088;
wire n10089;
wire n10090;
wire n10091;
wire n10092;
wire n10093;
wire n10094;
wire n10095;
wire n10096;
wire n10097;
wire n10098;
wire n10099;
wire n10100;
wire n10101;
wire n10102;
wire n10103;
wire n10104;
wire n10105;
wire n10106;
wire n10107;
wire n10108;
wire n10110;
wire n10111;
wire n10112;
wire n10113;
wire n10114;
wire n10115;
wire n10116;
wire n10117;
wire n10118;
wire n10119;
wire n10120;
wire n10121;
wire n10122;
wire n10123;
wire n10124;
wire n10125;
wire n10126;
wire n10127;
wire n10128;
wire n10129;
wire n10130;
wire n10131;
wire n10132;
wire n10133;
wire n10134;
wire n10135;
wire n10136;
wire n10137;
wire n10138;
wire n10139;
wire n10140;
wire n10141;
wire n10142;
wire n10143;
wire n10144;
wire n10145;
wire n10146;
wire n10147;
wire n10148;
wire n10149;
wire n10150;
wire n10151;
wire n10152;
wire n10153;
wire n10154;
wire n10155;
wire n10156;
wire n10157;
wire n10158;
wire n10159;
wire n10160;
wire n10161;
wire n10162;
wire n10163;
wire n10164;
wire n10165;
wire n10167;
wire n10168;
wire n10169;
wire n10170;
wire n10171;
wire n10172;
wire n10173;
wire n10174;
wire n10175;
wire n10176;
wire n10177;
wire n10178;
wire n10179;
wire n10180;
wire n10181;
wire n10182;
wire n10183;
wire n10184;
wire n10185;
wire n10186;
wire n10187;
wire n10188;
wire n10189;
wire n10190;
wire n10191;
wire n10192;
wire n10193;
wire n10194;
wire n10195;
wire n10196;
wire n10197;
wire n10198;
wire n10199;
wire n10200;
wire n10201;
wire n10202;
wire n10203;
wire n10204;
wire n10205;
wire n10206;
wire n10207;
wire n10208;
wire n10209;
wire n10210;
wire n10211;
wire n10212;
wire n10213;
wire n10214;
wire n10215;
wire n10216;
wire n10217;
wire n10218;
wire n10219;
wire n10221;
wire n10222;
wire n10223;
wire n10224;
wire n10225;
wire n10228;
wire n10229;
wire n10230;
wire n10231;
wire n10232;
wire n10233;
wire n10234;
wire n10235;
wire n10236;
wire n10237;
wire n10238;
wire n10239;
wire n10240;
wire n10241;
wire n10242;
wire n10243;
wire n10244;
wire n10245;
wire n10246;
wire n10247;
wire n10248;
wire n10249;
wire n10250;
wire n10251;
wire n10252;
wire n10253;
wire n10254;
wire n10255;
wire n10257;
wire n10258;
wire n10259;
wire n10260;
wire n10261;
wire n10262;
wire n10264;
wire n10265;
wire n10266;
wire n10267;
wire n10268;
wire n10269;
wire n10270;
wire n10271;
wire n10272;
wire n10273;
wire n10274;
wire n10275;
wire n10276;
wire n10277;
wire n10278;
wire n10279;
wire n10280;
wire n10281;
wire n10282;
wire n10283;
wire n10284;
wire n10285;
wire n10286;
wire n10287;
wire n10288;
wire n10289;
wire n10290;
wire n10291;
wire n10292;
wire n10293;
wire n10294;
wire n10295;
wire n10296;
wire n10297;
wire n10298;
wire n10299;
wire n10300;
wire n10301;
wire n10302;
wire n10303;
wire n10304;
wire n10305;
wire n10306;
wire n10307;
wire n10308;
wire n10309;
wire n10310;
wire n10311;
wire n10312;
wire n10315;
wire n10316;
wire n10317;
wire n10318;
wire n10319;
wire n10320;
wire n10321;
wire n10322;
wire n10323;
wire n10324;
wire n10325;
wire n10326;
wire n10327;
wire n10328;
wire n10329;
wire n10330;
wire n10331;
wire n10332;
wire n10333;
wire n10334;
wire n10335;
wire n10336;
wire n10337;
wire n10338;
wire n10339;
wire n10341;
wire n10342;
wire n10343;
wire n10344;
wire n10345;
wire n10346;
wire n10347;
wire n10348;
wire n10349;
wire n10350;
wire n10351;
wire n10352;
wire n10353;
wire n10354;
wire n10355;
wire n10356;
wire n10357;
wire n10358;
wire n10359;
wire n10360;
wire n10361;
wire n10362;
wire n10363;
wire n10364;
wire n10365;
wire n10366;
wire n10367;
wire n10368;
wire n10369;
wire n10370;
wire n10371;
wire n10372;
wire n10373;
wire n10374;
wire n10375;
wire n10376;
wire n10377;
wire n10378;
wire n10379;
wire n10380;
wire n10381;
wire n10382;
wire n10383;
wire n10384;
wire n10385;
wire n10386;
wire n10387;
wire n10388;
wire n10389;
wire n10390;
wire n10391;
wire n10392;
wire n10393;
wire n10394;
wire n10395;
wire n10396;
wire n10397;
wire n10398;
wire n10399;
wire n10400;
wire n10401;
wire n10402;
wire n10404;
wire n10405;
wire n10406;
wire n10407;
wire n10408;
wire n10409;
wire n10410;
wire n10411;
wire n10412;
wire n10414;
wire n10415;
wire n10416;
wire n10417;
wire n10418;
wire n10419;
wire n10420;
wire n10421;
wire n10422;
wire n10423;
wire n10424;
wire n10425;
wire n10426;
wire n10427;
wire n10428;
wire n10429;
wire n10430;
wire n10431;
wire n10432;
wire n10433;
wire n10434;
wire n10435;
wire n10436;
wire n10437;
wire n10438;
wire n10439;
wire n10440;
wire n10441;
wire n10442;
wire n10443;
wire n10444;
wire n10445;
wire n10446;
wire n10447;
wire n10448;
wire n10449;
wire n10450;
wire n10451;
wire n10452;
wire n10453;
wire n10454;
wire n10455;
wire n10456;
wire n10457;
wire n10458;
wire n10459;
wire n10460;
wire n10461;
wire n10462;
wire n10463;
wire n10464;
wire n10465;
wire n10466;
wire n10467;
wire n10468;
wire n10469;
wire n10470;
wire n10471;
wire n10472;
wire n10473;
wire n10474;
wire n10475;
wire n10476;
wire n10477;
wire n10478;
wire n10479;
wire n10480;
wire n10481;
wire n10482;
wire n10483;
wire n10484;
wire n10485;
wire n10486;
wire n10487;
wire n10488;
wire n10489;
wire n10490;
wire n10491;
wire n10492;
wire n10493;
wire n10494;
wire n10495;
wire n10496;
wire n10497;
wire n10498;
wire n10499;
wire n10500;
wire n10501;
wire n10502;
wire n10503;
wire n10504;
wire n10505;
wire n10506;
wire n10507;
wire n10508;
wire n10509;
wire n10510;
wire n10511;
wire n10512;
wire n10513;
wire n10514;
wire n10515;
wire n10516;
wire n10517;
wire n10518;
wire n10519;
wire n10520;
wire n10521;
wire n10522;
wire n10523;
wire n10524;
wire n10526;
wire n10527;
wire n10528;
wire n10529;
wire n10530;
wire n10531;
wire n10532;
wire n10533;
wire n10534;
wire n10535;
wire n10536;
wire n10537;
wire n10538;
wire n10539;
wire n10540;
wire n10541;
wire n10542;
wire n10543;
wire n10544;
wire n10545;
wire n10546;
wire n10547;
wire n10548;
wire n10549;
wire n10550;
wire n10551;
wire n10552;
wire n10553;
wire n10554;
wire n10555;
wire n10556;
wire n10557;
wire n10559;
wire n10560;
wire n10561;
wire n10562;
wire n10563;
wire n10564;
wire n10565;
wire n10566;
wire n10567;
wire n10568;
wire n10569;
wire n10570;
wire n10571;
wire n10572;
wire n10573;
wire n10574;
wire n10575;
wire n10576;
wire n10577;
wire n10578;
wire n10579;
wire n10580;
wire n10581;
wire n10582;
wire n10583;
wire n10584;
wire n10585;
wire n10586;
wire n10587;
wire n10588;
wire n10589;
wire n10590;
wire n10591;
wire n10592;
wire n10593;
wire n10594;
wire n10595;
wire n10596;
wire n10597;
wire n10598;
wire n10599;
wire n10600;
wire n10601;
wire n10602;
wire n10603;
wire n10604;
wire n10605;
wire n10606;
wire n10607;
wire n10608;
wire n10609;
wire n10610;
wire n10611;
wire n10612;
wire n10613;
wire n10614;
wire n10615;
wire n10616;
wire n10617;
wire n10618;
wire n10619;
wire n10620;
wire n10621;
wire n10622;
wire n10623;
wire n10624;
wire n10625;
wire n10626;
wire n10627;
wire n10628;
wire n10629;
wire n10630;
wire n10631;
wire n10632;
wire n10633;
wire n10634;
wire n10635;
wire n10636;
wire n10637;
wire n10638;
wire n10639;
wire n10640;
wire n10641;
wire n10642;
wire n10643;
wire n10644;
wire n10645;
wire n10646;
wire n10647;
wire n10648;
wire n10649;
wire n10650;
wire n10651;
wire n10652;
wire n10653;
wire n10654;
wire n10655;
wire n10656;
wire n10657;
wire n10658;
wire n10659;
wire n10660;
wire n10661;
wire n10662;
wire n10663;
wire n10664;
wire n10665;
wire n10666;
wire n10667;
wire n10668;
wire n10669;
wire n10670;
wire n10671;
wire n10672;
wire n10673;
wire n10674;
wire n10675;
wire n10676;
wire n10677;
wire n10678;
wire n10679;
wire n10680;
wire n10681;
wire n10682;
wire n10683;
wire n10684;
wire n10685;
wire n10686;
wire n10687;
wire n10688;
wire n10689;
wire n10690;
wire n10691;
wire n10692;
wire n10693;
wire n10694;
wire n10695;
wire n10696;
wire n10697;
wire n10698;
wire n10699;
wire n10700;
wire n10701;
wire n10702;
wire n10703;
wire n10704;
wire n10705;
wire n10706;
wire n10707;
wire n10708;
wire n10709;
wire n10710;
wire n10711;
wire n10712;
wire n10713;
wire n10714;
wire n10715;
wire n10716;
wire n10717;
wire n10718;
wire n10719;
wire n10720;
wire n10721;
wire n10722;
wire n10723;
wire n10724;
wire n10725;
wire n10726;
wire n10727;
wire n10728;
wire n10729;
wire n10730;
wire n10731;
wire n10732;
wire n10733;
wire n10734;
wire n10735;
wire n10736;
wire n10737;
wire n10738;
wire n10739;
wire n10740;
wire n10741;
wire n10742;
wire n10743;
wire n10744;
wire n10745;
wire n10746;
wire n10747;
wire n10748;
wire n10749;
wire n10750;
wire n10751;
wire n10752;
wire n10753;
wire n10754;
wire n10755;
wire n10756;
wire n10757;
wire n10758;
wire n10759;
wire n10760;
wire n10761;
wire n10762;
wire n10763;
wire n10764;
wire n10765;
wire n10766;
wire n10767;
wire n10768;
wire n10769;
wire n10770;
wire n10771;
wire n10772;
wire n10773;
wire n10774;
wire n10775;
wire n10776;
wire n10777;
wire n10778;
wire n10779;
wire n10780;
wire n10781;
wire n10782;
wire n10783;
wire n10784;
wire n10785;
wire n10786;
wire n10787;
wire n10788;
wire n10789;
wire n10790;
wire n10791;
wire n10792;
wire n10793;
wire n10794;
wire n10795;
wire n10796;
wire n10797;
wire n10798;
wire n10799;
wire n10800;
wire n10801;
wire n10802;
wire n10803;
wire n10804;
wire n10805;
wire n10806;
wire n10807;
wire n10808;
wire n10809;
wire n10810;
wire n10811;
wire n10812;
wire n10813;
wire n10814;
wire n10815;
wire n10816;
wire n10817;
wire n10818;
wire n10819;
wire n10820;
wire n10821;
wire n10822;
wire n10823;
wire n10824;
wire n10825;
wire n10826;
wire n10827;
wire n10828;
wire n10829;
wire n10830;
wire n10831;
wire n10832;
wire n10833;
wire n10834;
wire n10835;
wire n10836;
wire n10837;
wire n10838;
wire n10839;
wire n10840;
wire n10841;
wire n10842;
wire n10843;
wire n10844;
wire n10845;
wire n10846;
wire n10847;
wire n10848;
wire n10849;
wire n10850;
wire n10851;
wire n10852;
wire n10853;
wire n10854;
wire n10855;
wire n10856;
wire n10857;
wire n10858;
wire n10859;
wire n10860;
wire n10861;
wire n10862;
wire n10863;
wire n10864;
wire n10865;
wire n10866;
wire n10867;
wire n10868;
wire n10869;
wire n10870;
wire n10871;
wire n10872;
wire n10873;
wire n10874;
wire n10875;
wire n10876;
wire n10877;
wire n10878;
wire n10879;
wire n10880;
wire n10881;
wire n10882;
wire n10883;
wire n10884;
wire n10885;
wire n10886;
wire n10887;
wire n10888;
wire n10889;
wire n10890;
wire n10891;
wire n10892;
wire n10893;
wire n10894;
wire n10895;
wire n10896;
wire n10897;
wire n10898;
wire n10899;
wire n10900;
wire n10901;
wire n10902;
wire n10903;
wire n10904;
wire n10905;
wire n10906;
wire n10907;
wire n10908;
wire n10909;
wire n10910;
wire n10911;
wire n10912;
wire n10913;
wire n10914;
wire n10915;
wire n10916;
wire n10917;
wire n10918;
wire n10919;
wire n10920;
wire n10921;
wire n10922;
wire n10923;
wire n10924;
wire n10925;
wire n10926;
wire n10927;
wire n10928;
wire n10929;
wire n10930;
wire n10931;
wire n10932;
wire n10933;
wire n10934;
wire n10935;
wire n10936;
wire n10937;
wire n10938;
wire n10939;
wire n10940;
wire n10941;
wire n10942;
wire n10943;
wire n10944;
wire n10945;
wire n10946;
wire n10947;
wire n10948;
wire n10949;
wire n10950;
wire n10951;
wire n10952;
wire n10953;
wire n10954;
wire n10955;
wire n10956;
wire n10957;
wire n10958;
wire n10959;
wire n10960;
wire n10961;
wire n10962;
wire n10963;
wire n10964;
wire n10965;
wire n10966;
wire n10967;
wire n10968;
wire n10969;
wire n10970;
wire n10971;
wire n10972;
wire n10973;
wire n10974;
wire n10975;
wire n10976;
wire n10977;
wire n10978;
wire n10979;
wire n10980;
wire n10981;
wire n10982;
wire n10983;
wire n10984;
wire n10985;
wire n10986;
wire n10987;
wire n10988;
wire n10989;
wire n10990;
wire n10991;
wire n10992;
wire n10993;
wire n10994;
wire n10995;
wire n10996;
wire n10997;
wire n10998;
wire n10999;
wire n11000;
wire n11001;
wire n11002;
wire n11003;
wire n11004;
wire n11005;
wire n11006;
wire n11007;
wire n11008;
wire n11009;
wire n11010;
wire n11011;
wire n11012;
wire n11013;
wire n11014;
wire n11015;
wire n11016;
wire n11017;
wire n11018;
wire n11019;
wire n11020;
wire n11021;
wire n11022;
wire n11023;
wire n11024;
wire n11025;
wire n11026;
wire n11027;
wire n11028;
wire n11029;
wire n11030;
wire n11031;
wire n11032;
wire n11033;
wire n11034;
wire n11035;
wire n11036;
wire n11037;
wire n11038;
wire n11039;
wire n11040;
wire n11041;
wire n11042;
wire n11043;
wire n11044;
wire n11045;
wire n11046;
wire n11047;
wire n11048;
wire n11049;
wire n11050;
wire n11051;
wire n11052;
wire n11053;
wire n11054;
wire n11055;
wire n11056;
wire n11057;
wire n11058;
wire n11059;
wire n11060;
wire n11061;
wire n11062;
wire n11063;
wire n11064;
wire n11065;
wire n11066;
wire n11067;
wire n11068;
wire n11069;
wire n11070;
wire n11071;
wire n11072;
wire n11073;
wire n11074;
wire n11075;
wire n11076;
wire n11077;
wire n11078;
wire n11079;
wire n11080;
wire n11081;
wire n11082;
wire n11083;
wire n11084;
wire n11085;
wire n11086;
wire n11087;
wire n11088;
wire n11089;
wire n11090;
wire n11091;
wire n11092;
wire n11093;
wire n11094;
wire n11095;
wire n11096;
wire n11097;
wire n11098;
wire n11099;
wire n11100;
wire n11101;
wire n11102;
wire n11103;
wire n11104;
wire n11105;
wire n11106;
wire n11107;
wire n11108;
wire n11109;
wire n11110;
wire n11111;
wire n11112;
wire n11113;
wire n11114;
wire n11115;
wire n11116;
wire n11117;
wire n11118;
wire n11119;
wire n11120;
wire n11121;
wire n11122;
wire n11123;
wire n11124;
wire n11125;
wire n11126;
wire n11127;
wire n11128;
wire n11129;
wire n11130;
wire n11131;
wire n11132;
wire n11133;
wire n11134;
wire n11135;
wire n11136;
wire n11137;
wire n11138;
wire n11139;
wire n11140;
wire n11141;
wire n11142;
wire n11143;
wire n11144;
wire n11145;
wire n11146;
wire n11147;
wire n11148;
wire n11149;
wire n11150;
wire n11151;
wire n11152;
wire n11153;
wire n11154;
wire n11155;
wire n11156;
wire n11157;
wire n11158;
wire n11159;
wire n11160;
wire n11161;
wire n11162;
wire n11163;
wire n11164;
wire n11165;
wire n11166;
wire n11167;
wire n11168;
wire n11169;
wire n11170;
wire n11171;
wire n11172;
wire n11173;
wire n11174;
wire n11175;
wire n11176;
wire n11177;
wire n11178;
wire n11179;
wire n11180;
wire n11181;
wire n11182;
wire n11183;
wire n11184;
wire n11185;
wire n11186;
wire n11187;
wire n11188;
wire n11189;
wire n11190;
wire n11191;
wire n11192;
wire n11193;
wire n11194;
wire n11195;
wire n11196;
wire n11197;
wire n11198;
wire n11199;
wire n11200;
wire n11201;
wire n11202;
wire n11203;
wire n11204;
wire n11205;
wire n11206;
wire n11207;
wire n11208;
wire n11209;
wire n11210;
wire n11211;
wire n11212;
wire n11213;
wire n11214;
wire n11215;
wire n11216;
wire n11217;
wire n11218;
wire n11219;
wire n11220;
wire n11221;
wire n11222;
wire n11223;
wire n11224;
wire n11225;
wire n11226;
wire n11227;
wire n11228;
wire n11229;
wire n11230;
wire n11231;
wire n11232;
wire n11233;
wire n11234;
wire n11235;
wire n11236;
wire n11237;
wire n11238;
wire n11239;
wire n11241;
wire n11242;
wire n11243;
wire n11244;
wire n11245;
wire n11246;
wire n11247;
wire n11248;
wire n11249;
wire n11250;
wire n11251;
wire n11252;
wire n11253;
wire n11254;
wire n11255;
wire n11256;
wire n11257;
wire n11258;
wire n11259;
wire n11260;
wire n11261;
wire n11262;
wire n11263;
wire n11264;
wire n11265;
wire n11266;
wire n11267;
wire n11268;
wire n11269;
wire n11270;
wire n11271;
wire n11272;
wire n11273;
wire n11274;
wire n11275;
wire n11276;
wire n11277;
wire n11278;
wire n11279;
wire n11280;
wire n11281;
wire n11283;
wire n11284;
wire n11285;
wire n11286;
wire n11287;
wire n11288;
wire n11289;
wire n11290;
wire n11291;
wire n11292;
wire n11293;
wire n11294;
wire n11295;
wire n11296;
wire n11297;
wire n11298;
wire n11299;
wire n11300;
wire n11301;
wire n11302;
wire n11303;
wire n11304;
wire n11305;
wire n11306;
wire n11307;
wire n11308;
wire n11309;
wire n11310;
wire n11311;
wire n11312;
wire n11313;
wire n11314;
wire n11315;
wire n11316;
wire n11317;
wire n11318;
wire n11319;
wire n11320;
wire n11321;
wire n11322;
wire n11323;
wire n11324;
wire n11325;
wire n11326;
wire n11327;
wire n11328;
wire n11329;
wire n11330;
wire n11331;
wire n11332;
wire n11333;
wire n11334;
wire n11335;
wire n11336;
wire n11337;
wire n11338;
wire n11339;
wire n11340;
wire n11341;
wire n11342;
wire n11343;
wire n11344;
wire n11345;
wire n11346;
wire n11347;
wire n11348;
wire n11349;
wire n11350;
wire n11351;
wire n11352;
wire n11353;
wire n11354;
wire n11355;
wire n11356;
wire n11357;
wire n11358;
wire n11359;
wire n11360;
wire n11361;
wire n11362;
wire n11363;
wire n11364;
wire n11365;
wire n11366;
wire n11367;
wire n11368;
wire n11369;
wire n11370;
wire n11371;
wire n11372;
wire n11373;
wire n11374;
wire n11375;
wire n11376;
wire n11377;
wire n11378;
wire n11379;
wire n11380;
wire n11381;
wire n11382;
wire n11383;
wire n11384;
wire n11385;
wire n11386;
wire n11387;
wire n11388;
wire n11389;
wire n11390;
wire n11391;
wire n11392;
wire n11393;
wire n11394;
wire n11395;
wire n11396;
wire n11397;
wire n11398;
wire n11399;
wire n11400;
wire n11401;
wire n11402;
wire n11403;
wire n11404;
wire n11405;
wire n11406;
wire n11407;
wire n11408;
wire n11409;
wire n11410;
wire n11411;
wire n11412;
wire n11413;
wire n11414;
wire n11415;
wire n11416;
wire n11417;
wire n11418;
wire n11419;
wire n11420;
wire n11421;
wire n11422;
wire n11423;
wire n11424;
wire n11425;
wire n11426;
wire n11427;
wire n11428;
wire n11429;
wire n11430;
wire n11431;
wire n11432;
wire n11433;
wire n11434;
wire n11435;
wire n11436;
wire n11437;
wire n11438;
wire n11439;
wire n11440;
wire n11441;
wire n11442;
wire n11443;
wire n11444;
wire n11445;
wire n11446;
wire n11447;
wire n11448;
wire n11449;
wire n11450;
wire n11451;
wire n11452;
wire n11453;
wire n11454;
wire n11455;
wire n11456;
wire n11457;
wire n11458;
wire n11459;
wire n11460;
wire n11461;
wire n11462;
wire n11463;
wire n11464;
wire n11465;
wire n11466;
wire n11467;
wire n11468;
wire n11469;
wire n11470;
wire n11471;
wire n11472;
wire n11473;
wire n11474;
wire n11475;
wire n11476;
wire n11477;
wire n11478;
wire n11479;
wire n11480;
wire n11481;
wire n11482;
wire n11483;
wire n11484;
wire n11485;
wire n11486;
wire n11487;
wire n11488;
wire n11489;
wire n11490;
wire n11491;
wire n11492;
wire n11493;
wire n11494;
wire n11495;
wire n11496;
wire n11497;
wire n11498;
wire n11499;
wire n11500;
wire n11501;
wire n11502;
wire n11503;
wire n11504;
wire n11505;
wire n11506;
wire n11507;
wire n11508;
wire n11510;
wire n11511;
wire n11512;
wire n11513;
wire n11514;
wire n11515;
wire n11516;
wire n11517;
wire n11518;
wire n11519;
wire n11520;
wire n11521;
wire n11522;
wire n11523;
wire n11524;
wire n11525;
wire n11526;
wire n11527;
wire n11528;
wire n11529;
wire n11530;
wire n11531;
wire n11532;
wire n11533;
wire n11534;
wire n11535;
wire n11536;
wire n11537;
wire n11538;
wire n11539;
wire n11540;
wire n11541;
wire n11542;
wire n11543;
wire n11544;
wire n11545;
wire n11546;
wire n11547;
wire n11548;
wire n11549;
wire n11550;
wire n11551;
wire n11552;
wire n11553;
wire n11554;
wire n11555;
wire n11556;
wire n11557;
wire n11558;
wire n11559;
wire n11560;
wire n11561;
wire n11562;
wire n11564;
wire n11565;
wire n11566;
wire n11567;
wire n11569;
wire n11570;
wire n11571;
wire n11572;
wire n11573;
wire n11574;
wire n11575;
wire n11576;
wire n11577;
wire n11578;
wire n11579;
wire n11580;
wire n11581;
wire n11582;
wire n11583;
wire n11584;
wire n11585;
wire n11586;
wire n11587;
wire n11588;
wire n11589;
wire n11590;
wire n11591;
wire n11592;
wire n11593;
wire n11594;
wire n11595;
wire n11596;
wire n11597;
wire n11598;
wire n11600;
wire n11601;
wire n11602;
wire n11603;
wire n11604;
wire n11605;
wire n11606;
wire n11607;
wire n11608;
wire n11609;
wire n11610;
wire n11611;
wire n11612;
wire n11613;
wire n11614;
wire n11615;
wire n11616;
wire n11617;
wire n11618;
wire n11619;
wire n11620;
wire n11621;
wire n11622;
wire n11623;
wire n11624;
wire n11625;
wire n11626;
wire n11627;
wire n11628;
wire n11629;
wire n11630;
wire n11631;
wire n11632;
wire n11633;
wire n11634;
wire n11635;
wire n11636;
wire n11637;
wire n11638;
wire n11639;
wire n11640;
wire n11641;
wire n11642;
wire n11643;
wire n11644;
wire n11645;
wire n11646;
wire n11647;
wire n11648;
wire n11649;
wire n11650;
wire n11651;
wire n11652;
wire n11653;
wire n11654;
wire n11655;
wire n11656;
wire n11657;
wire n11658;
wire n11659;
wire n11660;
wire n11661;
wire n11662;
wire n11663;
wire n11664;
wire n11665;
wire n11666;
wire n11667;
wire n11668;
wire n11669;
wire n11670;
wire n11671;
wire n11672;
wire n11673;
wire n11674;
wire n11675;
wire n11676;
wire n11677;
wire n11678;
wire n11679;
wire n11680;
wire n11681;
wire n11682;
wire n11683;
wire n11684;
wire n11685;
wire n11686;
wire n11687;
wire n11688;
wire n11689;
wire n11690;
wire n11691;
wire n11692;
wire n11693;
wire n11694;
wire n11695;
wire n11696;
wire n11697;
wire n11698;
wire n11699;
wire n11700;
wire n11701;
wire n11702;
wire n11703;
wire n11704;
wire n11705;
wire n11706;
wire n11707;
wire n11708;
wire n11709;
wire n11710;
wire n11711;
wire n11712;
wire n11713;
wire n11714;
wire n11715;
wire n11716;
wire n11717;
wire n11718;
wire n11719;
wire n11720;
wire n11721;
wire n11722;
wire n11723;
wire n11724;
wire n11725;
wire n11726;
wire n11727;
wire n11728;
wire n11729;
wire n11730;
wire n11731;
wire n11732;
wire n11733;
wire n11734;
wire n11735;
wire n11736;
wire n11737;
wire n11738;
wire n11739;
wire n11740;
wire n11741;
wire n11742;
wire n11743;
wire n11744;
wire n11745;
wire n11746;
wire n11747;
wire n11748;
wire n11749;
wire n11750;
wire n11751;
wire n11752;
wire n11753;
wire n11754;
wire n11755;
wire n11756;
wire n11757;
wire n11758;
wire n11759;
wire n11760;
wire n11761;
wire n11762;
wire n11763;
wire n11764;
wire n11765;
wire n11766;
wire n11767;
wire n11768;
wire n11769;
wire n11770;
wire n11771;
wire n11772;
wire n11773;
wire n11774;
wire n11775;
wire n11776;
wire n11777;
wire n11778;
wire n11779;
wire n11780;
wire n11781;
wire n11782;
wire n11783;
wire n11784;
wire n11785;
wire n11786;
wire n11787;
wire n11788;
wire n11789;
wire n11790;
wire n11791;
wire n11792;
wire n11793;
wire n11794;
wire n11795;
wire n11796;
wire n11797;
wire n11798;
wire n11799;
wire n11800;
wire n11801;
wire n11802;
wire n11803;
wire n11804;
wire n11805;
wire n11806;
wire n11807;
wire n11808;
wire n11809;
wire n11810;
wire n11811;
wire n11812;
wire n11813;
wire n11814;
wire n11815;
wire n11816;
wire n11817;
wire n11818;
wire n11819;
wire n11820;
wire n11821;
wire n11822;
wire n11823;
wire n11824;
wire n11825;
wire n11826;
wire n11827;
wire n11828;
wire n11829;
wire n11830;
wire n11831;
wire n11832;
wire n11833;
wire n11834;
wire n11835;
wire n11836;
wire n11837;
wire n11838;
wire n11839;
wire n11840;
wire n11841;
wire n11842;
wire n11843;
wire n11844;
wire n11845;
wire n11846;
wire n11847;
wire n11848;
wire n11849;
wire n11850;
wire n11851;
wire n11852;
wire n11853;
wire n11854;
wire n11856;
wire n11857;
wire n11858;
wire n11859;
wire n11860;
wire n11861;
wire n11862;
wire n11863;
wire n11864;
wire n11865;
wire n11866;
wire n11867;
wire n11868;
wire n11869;
wire n11870;
wire n11871;
wire n11872;
wire n11873;
wire n11874;
wire n11875;
wire n11876;
wire n11877;
wire n11878;
wire n11879;
wire n11880;
wire n11881;
wire n11882;
wire n11883;
wire n11884;
wire n11885;
wire n11886;
wire n11887;
wire n11888;
wire n11889;
wire n11890;
wire n11891;
wire n11892;
wire n11893;
wire n11894;
wire n11895;
wire n11896;
wire n11897;
wire n11898;
wire n11899;
wire n11900;
wire n11901;
wire n11902;
wire n11903;
wire n11904;
wire n11905;
wire n11906;
wire n11907;
wire n11908;
wire n11909;
wire n11910;
wire n11911;
wire n11912;
wire n11913;
wire n11914;
wire n11915;
wire n11916;
wire n11917;
wire n11918;
wire n11919;
wire n11920;
wire n11921;
wire n11922;
wire n11923;
wire n11924;
wire n11925;
wire n11926;
wire n11927;
wire n11928;
wire n11929;
wire n11930;
wire n11931;
wire n11932;
wire n11933;
wire n11935;
wire n11936;
wire n11937;
wire n11938;
wire n11939;
wire n11940;
wire n11941;
wire n11942;
wire n11943;
wire n11944;
wire n11945;
wire n11946;
wire n11947;
wire n11948;
wire n11949;
wire n11950;
wire n11951;
wire n11952;
wire n11953;
wire n11954;
wire n11955;
wire n11956;
wire n11957;
wire n11958;
wire n11959;
wire n11960;
wire n11961;
wire n11962;
wire n11963;
wire n11964;
wire n11965;
wire n11966;
wire n11967;
wire n11968;
wire n11969;
wire n11970;
wire n11971;
wire n11972;
wire n11973;
wire n11974;
wire n11975;
wire n11976;
wire n11977;
wire n11978;
wire n11979;
wire n11980;
wire n11981;
wire n11982;
wire n11983;
wire n11984;
wire n11985;
wire n11986;
wire n11987;
wire n11988;
wire n11989;
wire n11990;
wire n11991;
wire n11992;
wire n11993;
wire n11994;
wire n11995;
wire n11996;
wire n11997;
wire n11998;
wire n11999;
wire n12000;
wire n12001;
wire n12002;
wire n12003;
wire n12004;
wire n12005;
wire n12006;
wire n12007;
wire n12008;
wire n12009;
wire n12010;
wire n12011;
wire n12012;
wire n12013;
wire n12014;
wire n12015;
wire n12016;
wire n12017;
wire n12018;
wire n12019;
wire n12020;
wire n12021;
wire n12022;
wire n12023;
wire n12024;
wire n12025;
wire n12026;
wire n12027;
wire n12028;
wire n12029;
wire n12030;
wire n12031;
wire n12032;
wire n12033;
wire n12034;
wire n12035;
wire n12036;
wire n12037;
wire n12038;
wire n12039;
wire n12040;
wire n12041;
wire n12042;
wire n12043;
wire n12044;
wire n12045;
wire n12046;
wire n12047;
wire n12048;
wire n12049;
wire n12050;
wire n12051;
wire n12052;
wire n12053;
wire n12054;
wire n12055;
wire n12056;
wire n12057;
wire n12058;
wire n12059;
wire n12060;
wire n12061;
wire n12062;
wire n12063;
wire n12065;
wire n12066;
wire n12067;
wire n12068;
wire n12069;
wire n12070;
wire n12071;
wire n12072;
wire n12073;
wire n12074;
wire n12075;
wire n12076;
wire n12077;
wire n12078;
wire n12079;
wire n12080;
wire n12081;
wire n12082;
wire n12083;
wire n12084;
wire n12085;
wire n12086;
wire n12087;
wire n12088;
wire n12089;
wire n12090;
wire n12091;
wire n12092;
wire n12093;
wire n12094;
wire n12095;
wire n12096;
wire n12097;
wire n12098;
wire n12099;
wire n12100;
wire n12101;
wire n12102;
wire n12103;
wire n12104;
wire n12105;
wire n12106;
wire n12107;
wire n12108;
wire n12109;
wire n12110;
wire n12111;
wire n12112;
wire n12113;
wire n12114;
wire n12115;
wire n12116;
wire n12117;
wire n12118;
wire n12119;
wire n12120;
wire n12121;
wire n12122;
wire n12123;
wire n12124;
wire n12125;
wire n12126;
wire n12127;
wire n12128;
wire n12129;
wire n12130;
wire n12131;
wire n12132;
wire n12133;
wire n12134;
wire n12135;
wire n12136;
wire n12137;
wire n12138;
wire n12139;
wire n12140;
wire n12141;
wire n12142;
wire n12143;
wire n12144;
wire n12145;
wire n12146;
wire n12147;
wire n12148;
wire n12149;
wire n12150;
wire n12151;
wire n12152;
wire n12153;
wire n12154;
wire n12155;
wire n12156;
wire n12157;
wire n12158;
wire n12159;
wire n12160;
wire n12161;
wire n12162;
wire n12163;
wire n12164;
wire n12165;
wire n12166;
wire n12167;
wire n12168;
wire n12169;
wire n12170;
wire n12171;
wire n12172;
wire n12173;
wire n12174;
wire n12175;
wire n12176;
wire n12177;
wire n12178;
wire n12179;
wire n12180;
wire n12181;
wire n12182;
wire n12183;
wire n12184;
wire n12185;
wire n12186;
wire n12187;
wire n12188;
wire n12189;
wire n12190;
wire n12191;
wire n12192;
wire n12193;
wire n12194;
wire n12195;
wire n12196;
wire n12197;
wire n12198;
wire n12199;
wire n12200;
wire n12201;
wire n12202;
wire n12203;
wire n12204;
wire n12205;
wire n12206;
wire n12207;
wire n12208;
wire n12211;
wire n12212;
wire n12213;
wire n12214;
wire n12215;
wire n12216;
wire n12217;
wire n12218;
wire n12219;
wire n12220;
wire n12221;
wire n12222;
wire n12223;
wire n12224;
wire n12225;
wire n12226;
wire n12227;
wire n12229;
wire n12230;
wire n12231;
wire n12232;
wire n12233;
wire n12234;
wire n12235;
wire n12236;
wire n12237;
wire n12238;
wire n12239;
wire n12240;
wire n12241;
wire n12242;
wire n12243;
wire n12244;
wire n12245;
wire n12246;
wire n12247;
wire n12248;
wire n12249;
wire n12250;
wire n12251;
wire n12252;
wire n12253;
wire n12254;
wire n12255;
wire n12256;
wire n12257;
wire n12258;
wire n12259;
wire n12260;
wire n12261;
wire n12262;
wire n12263;
wire n12264;
wire n12265;
wire n12266;
wire n12267;
wire n12268;
wire n12269;
wire n12270;
wire n12271;
wire n12272;
wire n12273;
wire n12274;
wire n12275;
wire n12276;
wire n12277;
wire n12278;
wire n12279;
wire n12280;
wire n12281;
wire n12282;
wire n12283;
wire n12284;
wire n12285;
wire n12286;
wire n12287;
wire n12288;
wire n12289;
wire n12290;
wire n12291;
wire n12292;
wire n12293;
wire n12294;
wire n12295;
wire n12296;
wire n12297;
wire n12298;
wire n12299;
wire n12300;
wire n12301;
wire n12302;
wire n12303;
wire n12304;
wire n12305;
wire n12306;
wire n12307;
wire n12308;
wire n12309;
wire n12310;
wire n12311;
wire n12312;
wire n12313;
wire n12314;
wire n12315;
wire n12316;
wire n12317;
wire n12318;
wire n12319;
wire n12320;
wire n12321;
wire n12322;
wire n12323;
wire n12324;
wire n12325;
wire n12326;
wire n12327;
wire n12328;
wire n12329;
wire n12330;
wire n12331;
wire n12332;
wire n12333;
wire n12334;
wire n12335;
wire n12336;
wire n12337;
wire n12338;
wire n12339;
wire n12340;
wire n12341;
wire n12342;
wire n12343;
wire n12344;
wire n12345;
wire n12346;
wire n12347;
wire n12348;
wire n12349;
wire n12350;
wire n12351;
wire n12352;
wire n12353;
wire n12354;
wire n12355;
wire n12356;
wire n12357;
wire n12358;
wire n12359;
wire n12360;
wire n12361;
wire n12362;
wire n12363;
wire n12364;
wire n12365;
wire n12366;
wire n12367;
wire n12368;
wire n12369;
wire n12370;
wire n12371;
wire n12372;
wire n12373;
wire n12374;
wire n12375;
wire n12376;
wire n12377;
wire n12378;
wire n12379;
wire n12380;
wire n12381;
wire n12382;
wire n12383;
wire n12384;
wire n12385;
wire n12386;
wire n12387;
wire n12388;
wire n12389;
wire n12390;
wire n12391;
wire n12392;
wire n12393;
wire n12394;
wire n12395;
wire n12396;
wire n12397;
wire n12398;
wire n12399;
wire n12400;
wire n12401;
wire n12402;
wire n12403;
wire n12404;
wire n12405;
wire n12406;
wire n12407;
wire n12408;
wire n12409;
wire n12410;
wire n12411;
wire n12412;
wire n12413;
wire n12414;
wire n12415;
wire n12416;
wire n12417;
wire n12418;
wire n12419;
wire n12420;
wire n12421;
wire n12422;
wire n12423;
wire n12424;
wire n12425;
wire n12426;
wire n12427;
wire n12428;
wire n12429;
wire n12430;
wire n12431;
wire n12432;
wire n12433;
wire n12434;
wire n12435;
wire n12436;
wire n12437;
wire n12438;
wire n12439;
wire n12440;
wire n12441;
wire n12442;
wire n12443;
wire n12444;
wire n12445;
wire n12446;
wire n12447;
wire n12448;
wire n12449;
wire n12450;
wire n12451;
wire n12452;
wire n12453;
wire n12454;
wire n12455;
wire n12456;
wire n12457;
wire n12458;
wire n12459;
wire n12460;
wire n12461;
wire n12462;
wire n12463;
wire n12464;
wire n12465;
wire n12466;
wire n12467;
wire n12468;
wire n12469;
wire n12470;
wire n12471;
wire n12472;
wire n12473;
wire n12474;
wire n12475;
wire n12476;
wire n12477;
wire n12478;
wire n12479;
wire n12480;
wire n12481;
wire n12482;
wire n12483;
wire n12484;
wire n12485;
wire n12486;
wire n12487;
wire n12488;
wire n12489;
wire n12490;
wire n12491;
wire n12492;
wire n12493;
wire n12494;
wire n12495;
wire n12496;
wire n12497;
wire n12498;
wire n12499;
wire n12500;
wire n12501;
wire n12502;
wire n12503;
wire n12504;
wire n12505;
wire n12506;
wire n12507;
wire n12508;
wire n12509;
wire n12510;
wire n12511;
wire n12512;
wire n12513;
wire n12514;
wire n12515;
wire n12516;
wire n12517;
wire n12518;
wire n12519;
wire n12520;
wire n12521;
wire n12522;
wire n12523;
wire n12524;
wire n12525;
wire n12526;
wire n12527;
wire n12528;
wire n12529;
wire n12530;
wire n12531;
wire n12532;
wire n12533;
wire n12534;
wire n12535;
wire n12536;
wire n12537;
wire n12538;
wire n12539;
wire n12540;
wire n12541;
wire n12542;
wire n12543;
wire n12544;
wire n12545;
wire n12546;
wire n12547;
wire n12548;
wire n12549;
wire n12550;
wire n12551;
wire n12552;
wire n12553;
wire n12554;
wire n12555;
wire n12556;
wire n12557;
wire n12558;
wire n12559;
wire n12560;
wire n12561;
wire n12562;
wire n12563;
wire n12564;
wire n12565;
wire n12566;
wire n12567;
wire n12568;
wire n12569;
wire n12570;
wire n12571;
wire n12572;
wire n12573;
wire n12574;
wire n12575;
wire n12576;
wire n12577;
wire n12578;
wire n12579;
wire n12580;
wire n12581;
wire n12582;
wire n12583;
wire n12584;
wire n12585;
wire n12586;
wire n12587;
wire n12588;
wire n12589;
wire n12590;
wire n12591;
wire n12592;
wire n12593;
wire n12594;
wire n12595;
wire n12596;
wire n12597;
wire n12598;
wire n12599;
wire n12600;
wire n12601;
wire n12602;
wire n12603;
wire n12604;
wire n12605;
wire n12606;
wire n12607;
wire n12608;
wire n12609;
wire n12610;
wire n12611;
wire n12612;
wire n12613;
wire n12614;
wire n12615;
wire n12616;
wire n12617;
wire n12618;
wire n12619;
wire n12620;
wire n12621;
wire n12622;
wire n12623;
wire n12624;
wire n12625;
wire n12626;
wire n12627;
wire n12628;
wire n12629;
wire n12630;
wire n12631;
wire n12632;
wire n12633;
wire n12634;
wire n12635;
wire n12636;
wire n12637;
wire n12638;
wire n12639;
wire n12640;
wire n12641;
wire n12642;
wire n12643;
wire n12644;
wire n12645;
wire n12646;
wire n12647;
wire n12648;
wire n12649;
wire n12650;
wire n12651;
wire n12652;
wire n12653;
wire n12654;
wire n12655;
wire n12656;
wire n12657;
wire n12658;
wire n12659;
wire n12660;
wire n12661;
wire n12662;
wire n12663;
wire n12664;
wire n12665;
wire n12666;
wire n12667;
wire n12668;
wire n12669;
wire n12670;
wire n12671;
wire n12672;
wire n12673;
wire n12674;
wire n12675;
wire n12676;
wire n12677;
wire n12678;
wire n12679;
wire n12680;
wire n12681;
wire n12682;
wire n12683;
wire n12684;
wire n12685;
wire n12686;
wire n12687;
wire n12688;
wire n12689;
wire n12690;
wire n12691;
wire n12692;
wire n12693;
wire n12694;
wire n12695;
wire n12696;
wire n12697;
wire n12698;
wire n12699;
wire n12700;
wire n12701;
wire n12702;
wire n12703;
wire n12704;
wire n12705;
wire n12706;
wire n12707;
wire n12708;
wire n12709;
wire n12710;
wire n12711;
wire n12712;
wire n12713;
wire n12714;
wire n12715;
wire n12716;
wire n12717;
wire n12718;
wire n12719;
wire n12720;
wire n12721;
wire n12722;
wire n12723;
wire n12724;
wire n12725;
wire n12726;
wire n12727;
wire n12728;
wire n12729;
wire n12730;
wire n12731;
wire n12732;
wire n12733;
wire n12734;
wire n12735;
wire n12736;
wire n12737;
wire n12738;
wire n12739;
wire n12740;
wire n12741;
wire n12742;
wire n12743;
wire n12744;
wire n12745;
wire n12746;
wire n12747;
wire n12748;
wire n12749;
wire n12750;
wire n12751;
wire n12752;
wire n12753;
wire n12754;
wire n12755;
wire n12756;
wire n12757;
wire n12758;
wire n12759;
wire n12760;
wire n12761;
wire n12763;
wire n12764;
wire n12765;
wire n12766;
wire n12767;
wire n12768;
wire n12769;
wire n12770;
wire n12771;
wire n12772;
wire n12773;
wire n12774;
wire n12775;
wire n12776;
wire n12777;
wire n12778;
wire n12779;
wire n12780;
wire n12781;
wire n12782;
wire n12783;
wire n12784;
wire n12785;
wire n12786;
wire n12787;
wire n12788;
wire n12789;
wire n12790;
wire n12791;
wire n12792;
wire n12793;
wire n12794;
wire n12795;
wire n12796;
wire n12797;
wire n12798;
wire n12799;
wire n12800;
wire n12801;
wire n12802;
wire n12803;
wire n12804;
wire n12805;
wire n12806;
wire n12807;
wire n12808;
wire n12809;
wire n12810;
wire n12811;
wire n12812;
wire n12813;
wire n12814;
wire n12815;
wire n12816;
wire n12817;
wire n12818;
wire n12819;
wire n12820;
wire n12821;
wire n12822;
wire n12823;
wire n12824;
wire n12825;
wire n12826;
wire n12827;
wire n12828;
wire n12829;
wire n12830;
wire n12831;
wire n12832;
wire n12833;
wire n12834;
wire n12835;
wire n12836;
wire n12837;
wire n12838;
wire n12839;
wire n12840;
wire n12841;
wire n12842;
wire n12843;
wire n12844;
wire n12845;
wire n12846;
wire n12847;
wire n12848;
wire n12849;
wire n12850;
wire n12851;
wire n12852;
wire n12853;
wire n12854;
wire n12855;
wire n12856;
wire n12857;
wire n12858;
wire n12859;
wire n12860;
wire n12861;
wire n12862;
wire n12863;
wire n12864;
wire n12865;
wire n12866;
wire n12867;
wire n12868;
wire n12869;
wire n12870;
wire n12871;
wire n12872;
wire n12873;
wire n12874;
wire n12875;
wire n12876;
wire n12877;
wire n12878;
wire n12879;
wire n12880;
wire n12881;
wire n12882;
wire n12883;
wire n12884;
wire n12885;
wire n12886;
wire n12887;
wire n12888;
wire n12889;
wire n12890;
wire n12891;
wire n12892;
wire n12893;
wire n12894;
wire n12895;
wire n12896;
wire n12897;
wire n12898;
wire n12899;
wire n12900;
wire n12901;
wire n12902;
wire n12903;
wire n12904;
wire n12905;
wire n12906;
wire n12907;
wire n12908;
wire n12909;
wire n12910;
wire n12911;
wire n12912;
wire n12913;
wire n12914;
wire n12915;
wire n12916;
wire n12917;
wire n12918;
wire n12919;
wire n12920;
wire n12921;
wire n12922;
wire n12923;
wire n12924;
wire n12925;
wire n12926;
wire n12927;
wire n12928;
wire n12929;
wire n12930;
wire n12931;
wire n12932;
wire n12933;
wire n12934;
wire n12935;
wire n12936;
wire n12937;
wire n12938;
wire n12939;
wire n12940;
wire n12941;
wire n12942;
wire n12943;
wire n12944;
wire n12945;
wire n12946;
wire n12947;
wire n12948;
wire n12949;
wire n12950;
wire n12951;
wire n12952;
wire n12953;
wire n12954;
wire n12955;
wire n12956;
wire n12957;
wire n12958;
wire n12959;
wire n12960;
wire n12961;
wire n12962;
wire n12963;
wire n12964;
wire n12965;
wire n12966;
wire n12967;
wire n12968;
wire n12969;
wire n12970;
wire n12971;
wire n12972;
wire n12973;
wire n12974;
wire n12975;
wire n12976;
wire n12977;
wire n12978;
wire n12979;
wire n12980;
wire n12981;
wire n12982;
wire n12983;
wire n12984;
wire n12985;
wire n12986;
wire n12987;
wire n12988;
wire n12989;
wire n12990;
wire n12991;
wire n12992;
wire n12993;
wire n12994;
wire n12995;
wire n12996;
wire n12997;
wire n12998;
wire n12999;
wire n13000;
wire n13001;
wire n13002;
wire n13003;
wire n13004;
wire n13005;
wire n13006;
wire n13007;
wire n13008;
wire n13009;
wire n13010;
wire n13011;
wire n13012;
wire n13013;
wire n13014;
wire n13015;
wire n13016;
wire n13017;
wire n13018;
wire n13019;
wire n13020;
wire n13021;
wire n13022;
wire n13023;
wire n13024;
wire n13025;
wire n13026;
wire n13027;
wire n13028;
wire n13029;
wire n13030;
wire n13031;
wire n13032;
wire n13033;
wire n13034;
wire n13035;
wire n13036;
wire n13037;
wire n13038;
wire n13039;
wire n13040;
wire n13041;
wire n13042;
wire n13043;
wire n13044;
wire n13045;
wire n13046;
wire n13047;
wire n13048;
wire n13049;
wire n13050;
wire n13051;
wire n13052;
wire n13053;
wire n13054;
wire n13055;
wire n13056;
wire n13057;
wire n13058;
wire n13059;
wire n13060;
wire n13061;
wire n13062;
wire n13063;
wire n13064;
wire n13065;
wire n13066;
wire n13067;
wire n13068;
wire n13069;
wire n13070;
wire n13071;
wire n13072;
wire n13073;
wire n13074;
wire n13075;
wire n13076;
wire n13077;
wire n13078;
wire n13079;
wire n13080;
wire n13081;
wire n13082;
wire n13083;
wire n13084;
wire n13085;
wire n13086;
wire n13087;
wire n13088;
wire n13089;
wire n13090;
wire n13091;
wire n13092;
wire n13093;
wire n13094;
wire n13095;
wire n13096;
wire n13097;
wire n13098;
wire n13099;
wire n13100;
wire n13101;
wire n13102;
wire n13103;
wire n13104;
wire n13105;
wire n13106;
wire n13107;
wire n13108;
wire n13109;
wire n13110;
wire n13111;
wire n13112;
wire n13113;
wire n13114;
wire n13115;
wire n13116;
wire n13117;
wire n13118;
wire n13119;
wire n13120;
wire n13121;
wire n13122;
wire n13123;
wire n13124;
wire n13125;
wire n13126;
wire n13127;
wire n13128;
wire n13129;
wire n13130;
wire n13131;
wire n13132;
wire n13133;
wire n13134;
wire n13135;
wire n13136;
wire n13138;
wire n13139;
wire n13140;
wire n13141;
wire n13142;
wire n13143;
wire n13144;
wire n13145;
wire n13146;
wire n13147;
wire n13148;
wire n13149;
wire n13150;
wire n13151;
wire n13152;
wire n13153;
wire n13154;
wire n13155;
wire n13156;
wire n13157;
wire n13158;
wire n13159;
wire n13160;
wire n13161;
wire n13162;
wire n13163;
wire n13164;
wire n13165;
wire n13166;
wire n13167;
wire n13168;
wire n13169;
wire n13170;
wire n13171;
wire n13172;
wire n13173;
wire n13174;
wire n13175;
wire n13176;
wire n13177;
wire n13178;
wire n13179;
wire n13180;
wire n13181;
wire n13182;
wire n13183;
wire n13184;
wire n13185;
wire n13186;
wire n13187;
wire n13188;
wire n13189;
wire n13190;
wire n13191;
wire n13192;
wire n13193;
wire n13194;
wire n13195;
wire n13196;
wire n13197;
wire n13198;
wire n13199;
wire n13200;
wire n13201;
wire n13202;
wire n13203;
wire n13204;
wire n13205;
wire n13206;
wire n13207;
wire n13208;
wire n13209;
wire n13210;
wire n13211;
wire n13212;
wire n13213;
wire n13214;
wire n13215;
wire n13216;
wire n13217;
wire n13218;
wire n13219;
wire n13220;
wire n13221;
wire n13222;
wire n13223;
wire n13224;
wire n13225;
wire n13226;
wire n13227;
wire n13228;
wire n13229;
wire n13230;
wire n13231;
wire n13232;
wire n13233;
wire n13234;
wire n13235;
wire n13236;
wire n13237;
wire n13238;
wire n13239;
wire n13240;
wire n13241;
wire n13242;
wire n13243;
wire n13244;
wire n13245;
wire n13246;
wire n13247;
wire n13248;
wire n13249;
wire n13250;
wire n13251;
wire n13252;
wire n13253;
wire n13254;
wire n13255;
wire n13256;
wire n13257;
wire n13258;
wire n13259;
wire n13260;
wire n13261;
wire n13262;
wire n13263;
wire n13264;
wire n13265;
wire n13266;
wire n13267;
wire n13268;
wire n13269;
wire n13270;
wire n13271;
wire n13272;
wire n13273;
wire n13274;
wire n13275;
wire n13276;
wire n13277;
wire n13278;
wire n13279;
wire n13280;
wire n13281;
wire n13282;
wire n13283;
wire n13284;
wire n13285;
wire n13286;
wire n13287;
wire n13288;
wire n13289;
wire n13290;
wire n13291;
wire n13292;
wire n13293;
wire n13294;
wire n13295;
wire n13296;
wire n13297;
wire n13298;
wire n13299;
wire n13300;
wire n13301;
wire n13302;
wire n13303;
wire n13304;
wire n13305;
wire n13306;
wire n13307;
wire n13308;
wire n13309;
wire n13310;
wire n13311;
wire n13312;
wire n13313;
wire n13314;
wire n13315;
wire n13316;
wire n13317;
wire n13318;
wire n13319;
wire n13320;
wire n13321;
wire n13322;
wire n13323;
wire n13324;
wire n13325;
wire n13326;
wire n13327;
wire n13328;
wire n13329;
wire n13330;
wire n13331;
wire n13332;
wire n13333;
wire n13334;
wire n13335;
wire n13336;
wire n13337;
wire n13338;
wire n13339;
wire n13340;
wire n13341;
wire n13342;
wire n13343;
wire n13344;
wire n13345;
wire n13346;
wire n13347;
wire n13348;
wire n13349;
wire n13350;
wire n13351;
wire n13352;
wire n13353;
wire n13354;
wire n13355;
wire n13356;
wire n13357;
wire n13358;
wire n13359;
wire n13360;
wire n13361;
wire n13362;
wire n13363;
wire n13364;
wire n13365;
wire n13366;
wire n13367;
wire n13368;
wire n13369;
wire n13370;
wire n13371;
wire n13372;
wire n13373;
wire n13374;
wire n13375;
wire n13376;
wire n13377;
wire n13378;
wire n13379;
wire n13380;
wire n13381;
wire n13382;
wire n13383;
wire n13384;
wire n13385;
wire n13386;
wire n13387;
wire n13388;
wire n13389;
wire n13390;
wire n13391;
wire n13392;
wire n13393;
wire n13394;
wire n13395;
wire n13396;
wire n13397;
wire n13398;
wire n13399;
wire n13400;
wire n13401;
wire n13402;
wire n13403;
wire n13404;
wire n13405;
wire n13406;
wire n13407;
wire n13408;
wire n13409;
wire n13410;
wire n13411;
wire n13412;
wire n13413;
wire n13414;
wire n13415;
wire n13416;
wire n13417;
wire n13418;
wire n13419;
wire n13420;
wire n13421;
wire n13422;
wire n13423;
wire n13424;
wire n13425;
wire n13426;
wire n13427;
wire n13428;
wire n13429;
wire n13430;
wire n13431;
wire n13432;
wire n13433;
wire n13434;
wire n13435;
wire n13436;
wire n13437;
wire n13438;
wire n13439;
wire n13440;
wire n13441;
wire n13442;
wire n13443;
wire n13444;
wire n13445;
wire n13446;
wire n13447;
wire n13448;
wire n13449;
wire n13450;
wire n13451;
wire n13452;
wire n13453;
wire n13454;
wire n13455;
wire n13456;
wire n13457;
wire n13458;
wire n13459;
wire n13460;
wire n13461;
wire n13462;
wire n13463;
wire n13464;
wire n13465;
wire n13466;
wire n13467;
wire n13468;
wire n13469;
wire n13470;
wire n13471;
wire n13472;
wire n13473;
wire n13474;
wire n13475;
wire n13476;
wire n13477;
wire n13478;
wire n13479;
wire n13480;
wire n13481;
wire n13482;
wire n13483;
wire n13484;
wire n13485;
wire n13486;
wire n13487;
wire n13488;
wire n13489;
wire n13490;
wire n13491;
wire n13492;
wire n13493;
wire n13494;
wire n13495;
wire n13496;
wire n13497;
wire n13498;
wire n13499;
wire n13500;
wire n13501;
wire n13502;
wire n13503;
wire n13504;
wire n13505;
wire n13506;
wire n13507;
wire n13508;
wire n13509;
wire n13510;
wire n13511;
wire n13512;
wire n13513;
wire n13514;
wire n13515;
wire n13516;
wire n13517;
wire n13518;
wire n13519;
wire n13520;
wire n13521;
wire n13522;
wire n13523;
wire n13524;
wire n13525;
wire n13526;
wire n13527;
wire n13528;
wire n13529;
wire n13530;
wire n13531;
wire n13532;
wire n13533;
wire n13534;
wire n13535;
wire n13536;
wire n13537;
wire n13538;
wire n13539;
wire n13540;
wire n13541;
wire n13542;
wire n13543;
wire n13544;
wire n13545;
wire n13546;
wire n13547;
wire n13548;
wire n13549;
wire n13550;
wire n13551;
wire n13552;
wire n13553;
wire n13554;
wire n13555;
wire n13556;
wire n13557;
wire n13558;
wire n13559;
wire n13560;
wire n13561;
wire n13562;
wire n13563;
wire n13564;
wire n13565;
wire n13566;
wire n13567;
wire n13568;
wire n13569;
wire n13570;
wire n13571;
wire n13572;
wire n13573;
wire n13574;
wire n13575;
wire n13576;
wire n13577;
wire n13578;
wire n13579;
wire n13580;
wire n13581;
wire n13582;
wire n13583;
wire n13584;
wire n13585;
wire n13586;
wire n13587;
wire n13588;
wire n13589;
wire n13590;
wire n13591;
wire n13592;
wire n13593;
wire n13594;
wire n13595;
wire n13596;
wire n13597;
wire n13598;
wire n13599;
wire n13600;
wire n13601;
wire n13602;
wire n13603;
wire n13604;
wire n13605;
wire n13606;
wire n13607;
wire n13608;
wire n13609;
wire n13610;
wire n13611;
wire n13612;
wire n13613;
wire n13614;
wire n13615;
wire n13616;
wire n13617;
wire n13618;
wire n13619;
wire n13620;
wire n13621;
wire n13622;
wire n13623;
wire n13624;
wire n13625;
wire n13626;
wire n13627;
wire n13628;
wire n13629;
wire n13630;
wire n13631;
wire n13632;
wire n13633;
wire n13634;
wire n13635;
wire n13636;
wire n13637;
wire n13638;
wire n13639;
wire n13640;
wire n13641;
wire n13642;
wire n13643;
wire n13644;
wire n13645;
wire n13646;
wire n13647;
wire n13648;
wire n13649;
wire n13650;
wire n13651;
wire n13652;
wire n13653;
wire n13654;
wire n13655;
wire n13656;
wire n13657;
wire n13658;
wire n13659;
wire n13660;
wire n13661;
wire n13662;
wire n13663;
wire n13664;
wire n13665;
wire n13666;
wire n13667;
wire n13668;
wire n13669;
wire n13670;
wire n13671;
wire n13672;
wire n13673;
wire n13674;
wire n13675;
wire n13676;
wire n13677;
wire n13678;
wire n13679;
wire n13680;
wire n13681;
wire n13682;
wire n13683;
wire n13684;
wire n13685;
wire n13686;
wire n13687;
wire n13688;
wire n13689;
wire n13690;
wire n13691;
wire n13692;
wire n13693;
wire n13694;
wire n13695;
wire n13696;
wire n13697;
wire n13698;
wire n13699;
wire n13700;
wire n13701;
wire n13702;
wire n13703;
wire n13704;
wire n13705;
wire n13706;
wire n13707;
wire n13708;
wire n13709;
wire n13710;
wire n13711;
wire n13712;
wire n13713;
wire n13714;
wire n13715;
wire n13716;
wire n13717;
wire n13718;
wire n13719;
wire n13720;
wire n13721;
wire n13722;
wire n13723;
wire n13724;
wire n13725;
wire n13726;
wire n13727;
wire n13728;
wire n13729;
wire n13730;
wire n13731;
wire n13732;
wire n13733;
wire n13734;
wire n13735;
wire n13736;
wire n13737;
wire n13738;
wire n13739;
wire n13740;
wire n13741;
wire n13742;
wire n13743;
wire n13744;
wire n13745;
wire n13746;
wire n13747;
wire n13748;
wire n13749;
wire n13750;
wire n13751;
wire n13752;
wire n13753;
wire n13754;
wire n13755;
wire n13756;
wire n13757;
wire n13758;
wire n13759;
wire n13760;
wire n13761;
wire n13762;
wire n13763;
wire n13764;
wire n13765;
wire n13766;
wire n13767;
wire n13768;
wire n13769;
wire n13770;
wire n13771;
wire n13772;
wire n13773;
wire n13774;
wire n13775;
wire n13776;
wire n13777;
wire n13778;
wire n13779;
wire n13780;
wire n13781;
wire n13782;
wire n13783;
wire n13784;
wire n13785;
wire n13786;
wire n13787;
wire n13788;
wire n13789;
wire n13790;
wire n13791;
wire n13792;
wire n13793;
wire n13794;
wire n13795;
wire n13796;
wire n13797;
wire n13798;
wire n13799;
wire n13800;
wire n13801;
wire n13802;
wire n13803;
wire n13804;
wire n13805;
wire n13806;
wire n13807;
wire n13808;
wire n13809;
wire n13810;
wire n13811;
wire n13812;
wire n13813;
wire n13814;
wire n13815;
wire n13816;
wire n13817;
wire n13818;
wire n13819;
wire n13820;
wire n13821;
wire n13822;
wire n13823;
wire n13824;
wire n13825;
wire n13826;
wire n13827;
wire n13828;
wire n13829;
wire n13830;
wire n13831;
wire n13832;
wire n13833;
wire n13834;
wire n13835;
wire n13836;
wire n13837;
wire n13838;
wire n13839;
wire n13840;
wire n13841;
wire n13842;
wire n13843;
wire n13844;
wire n13845;
wire n13846;
wire n13847;
wire n13848;
wire n13849;
wire n13850;
wire n13851;
wire n13852;
wire n13853;
wire n13854;
wire n13855;
wire n13856;
wire n13857;
wire n13858;
wire n13859;
wire n13860;
wire n13861;
wire n13862;
wire n13863;
wire n13864;
wire n13865;
wire n13866;
wire n13867;
wire n13868;
wire n13869;
wire n13870;
wire n13871;
wire n13872;
wire n13873;
wire n13874;
wire n13875;
wire n13876;
wire n13877;
wire n13878;
wire n13879;
wire n13880;
wire n13881;
wire n13882;
wire n13883;
wire n13884;
wire n13885;
wire n13886;
wire n13887;
wire n13888;
wire n13889;
wire n13890;
wire n13891;
wire n13892;
wire n13893;
wire n13894;
wire n13895;
wire n13896;
wire n13897;
wire n13898;
wire n13899;
wire n13900;
wire n13901;
wire n13902;
wire n13903;
wire n13904;
wire n13905;
wire n13906;
wire n13907;
wire n13908;
wire n13909;
wire n13910;
wire n13911;
wire n13912;
wire n13913;
wire n13914;
wire n13915;
wire n13916;
wire n13917;
wire n13918;
wire n13919;
wire n13920;
wire n13921;
wire n13922;
wire n13923;
wire n13924;
wire n13925;
wire n13926;
wire n13927;
wire n13928;
wire n13929;
wire n13930;
wire n13931;
wire n13932;
wire n13933;
wire n13934;
wire n13935;
wire n13936;
wire n13937;
wire n13938;
wire n13939;
wire n13940;
wire n13941;
wire n13942;
wire n13943;
wire n13944;
wire n13945;
wire n13946;
wire n13947;
wire n13948;
wire n13949;
wire n13950;
wire n13951;
wire n13952;
wire n13953;
wire n13954;
wire n13955;
wire n13956;
wire n13957;
wire n13958;
wire n13959;
wire n13960;
wire n13961;
wire n13962;
wire n13963;
wire n13964;
wire n13965;
wire n13966;
wire n13967;
wire n13968;
wire n13969;
wire n13970;
wire n13971;
wire n13972;
wire n13973;
wire n13974;
wire n13975;
wire n13976;
wire n13977;
wire n13978;
wire n13979;
wire n13980;
wire n13981;
wire n13982;
wire n13983;
wire n13984;
wire n13985;
wire n13986;
wire n13987;
wire n13988;
wire n13989;
wire n13990;
wire n13991;
wire n13992;
wire n13993;
wire n13994;
wire n13995;
wire n13996;
wire n13997;
wire n13998;
wire n13999;
wire n14000;
wire n14001;
wire n14002;
wire n14003;
wire n14004;
wire n14005;
wire n14006;
wire n14007;
wire n14008;
wire n14009;
wire n14010;
wire n14011;
wire n14012;
wire n14013;
wire n14014;
wire n14015;
wire n14016;
wire n14017;
wire n14018;
wire n14019;
wire n14020;
wire n14021;
wire n14022;
wire n14023;
wire n14024;
wire n14025;
wire n14026;
wire n14027;
wire n14028;
wire n14029;
wire n14030;
wire n14031;
wire n14032;
wire n14033;
wire n14034;
wire n14035;
wire n14036;
wire n14037;
wire n14038;
wire n14039;
wire n14040;
wire n14041;
wire n14042;
wire n14043;
wire n14044;
wire n14045;
wire n14046;
wire n14047;
wire n14048;
wire n14049;
wire n14050;
wire n14051;
wire n14052;
wire n14053;
wire n14054;
wire n14055;
wire n14056;
wire n14057;
wire n14058;
wire n14059;
wire n14060;
wire n14061;
wire n14062;
wire n14063;
wire n14064;
wire n14065;
wire n14066;
wire n14067;
wire n14068;
wire n14069;
wire n14070;
wire n14071;
wire n14072;
wire n14073;
wire n14074;
wire n14075;
wire n14076;
wire n14077;
wire n14078;
wire n14079;
wire n14080;
wire n14081;
wire n14082;
wire n14083;
wire n14084;
wire n14085;
wire n14086;
wire n14087;
wire n14088;
wire n14089;
wire n14090;
wire n14091;
wire n14092;
wire n14093;
wire n14094;
wire n14095;
wire n14096;
wire n14097;
wire n14098;
wire n14099;
wire n14100;
wire n14101;
wire n14102;
wire n14103;
wire n14104;
wire n14105;
wire n14106;
wire n14107;
wire n14108;
wire n14109;
wire n14110;
wire n14111;
wire n14112;
wire n14113;
wire n14114;
wire n14115;
wire n14116;
wire n14117;
wire n14118;
wire n14119;
wire n14120;
wire n14121;
wire n14122;
wire n14123;
wire n14124;
wire n14125;
wire n14126;
wire n14127;
wire n14128;
wire n14129;
wire n14130;
wire n14131;
wire n14132;
wire n14133;
wire n14134;
wire n14135;
wire n14136;
wire n14137;
wire n14138;
wire n14139;
wire n14140;
wire n14141;
wire n14142;
wire n14143;
wire n14144;
wire n14145;
wire n14146;
wire n14147;
wire n14148;
wire n14149;
wire n14150;
wire n14151;
wire n14152;
wire n14153;
wire n14154;
wire n14155;
wire n14156;
wire n14157;
wire n14158;
wire n14159;
wire n14160;
wire n14161;
wire n14162;
wire n14163;
wire n14164;
wire n14165;
wire n14166;
wire n14167;
wire n14168;
wire n14169;
wire n14170;
wire n14171;
wire n14172;
wire n14173;
wire n14174;
wire n14175;
wire n14176;
wire n14177;
wire n14178;
wire n14179;
wire n14180;
wire n14181;
wire n14182;
wire n14183;
wire n14184;
wire n14185;
wire n14186;
wire n14187;
wire n14188;
wire n14189;
wire n14190;
wire n14191;
wire n14192;
wire n14193;
wire n14194;
wire n14195;
wire n14196;
wire n14197;
wire n14198;
wire n14199;
wire n14200;
wire n14201;
wire n14202;
wire n14203;
wire n14204;
wire n14205;
wire n14206;
wire n14207;
wire n14208;
wire n14209;
wire n14210;
wire n14211;
wire n14212;
wire n14213;
wire n14214;
wire n14215;
wire n14216;
wire n14217;
wire n14218;
wire n14219;
wire n14220;
wire n14221;
wire n14222;
wire n14223;
wire n14224;
wire n14225;
wire n14226;
wire n14227;
wire n14228;
wire n14229;
wire n14230;
wire n14231;
wire n14232;
wire n14233;
wire n14234;
wire n14235;
wire n14236;
wire n14237;
wire n14238;
wire n14239;
wire n14240;
wire n14241;
wire n14242;
wire n14243;
wire n14244;
wire n14245;
wire n14246;
wire n14247;
wire n14248;
wire n14249;
wire n14250;
wire n14251;
wire n14252;
wire n14253;
wire n14254;
wire n14255;
wire n14256;
wire n14257;
wire n14258;
wire n14259;
wire n14260;
wire n14261;
wire n14262;
wire n14263;
wire n14264;
wire n14265;
wire n14266;
wire n14267;
wire n14268;
wire n14269;
wire n14270;
wire n14271;
wire n14272;
wire n14273;
wire n14274;
wire n14275;
wire n14276;
wire n14277;
wire n14278;
wire n14279;
wire n14280;
wire n14281;
wire n14282;
wire n14283;
wire n14284;
wire n14285;
wire n14286;
wire n14287;
wire n14288;
wire n14289;
wire n14290;
wire n14291;
wire n14292;
wire n14293;
wire n14294;
wire n14295;
wire n14296;
wire n14297;
wire n14298;
wire n14299;
wire n14300;
wire n14301;
wire n14302;
wire n14303;
wire n14304;
wire n14305;
wire n14306;
wire n14307;
wire n14308;
wire n14309;
wire n14310;
wire n14311;
wire n14312;
wire n14313;
wire n14314;
wire n14315;
wire n14316;
wire n14317;
wire n14318;
wire n14319;
wire n14320;
wire n14321;
wire n14322;
wire n14323;
wire n14324;
wire n14325;
wire n14326;
wire n14327;
wire n14328;
wire n14329;
wire n14330;
wire n14331;
wire n14332;
wire n14333;
wire n14334;
wire n14335;
wire n14336;
wire n14337;
wire n14338;
wire n14339;
wire n14340;
wire n14341;
wire n14342;
wire n14343;
wire n14344;
wire n14345;
wire n14346;
wire n14347;
wire n14348;
wire n14349;
wire n14350;
wire n14351;
wire n14352;
wire n14353;
wire n14354;
wire n14355;
wire n14356;
wire n14357;
wire n14358;
wire n14359;
wire n14360;
wire n14361;
wire n14362;
wire n14363;
wire n14364;
wire n14365;
wire n14366;
wire n14367;
wire n14368;
wire n14369;
wire n14370;
wire n14371;
wire n14372;
wire n14373;
wire n14374;
wire n14375;
wire n14376;
wire n14377;
wire n14378;
wire n14379;
wire n14380;
wire n14381;
wire n14382;
wire n14383;
wire n14384;
wire n14385;
wire n14386;
wire n14387;
wire n14388;
wire n14389;
wire n14390;
wire n14391;
wire n14392;
wire n14393;
wire n14394;
wire n14395;
wire n14396;
wire n14397;
wire n14398;
wire n14399;
wire n14400;
wire n14401;
wire n14402;
wire n14403;
wire n14404;
wire n14405;
wire n14406;
wire n14407;
wire n14408;
wire n14409;
wire n14410;
wire n14411;
wire n14412;
wire n14413;
wire n14414;
wire n14415;
wire n14416;
wire n14417;
wire n14418;
wire n14419;
wire n14420;
wire n14421;
wire n14422;
wire n14423;
wire n14424;
wire n14425;
wire n14426;
wire n14427;
wire n14428;
wire n14429;
wire n14430;
wire n14431;
wire n14432;
wire n14433;
wire n14434;
wire n14435;
wire n14436;
wire n14437;
wire n14438;
wire n14439;
wire n14440;
wire n14441;
wire n14442;
wire n14443;
wire n14444;
wire n14445;
wire n14446;
wire n14447;
wire n14448;
wire n14449;
wire n14450;
wire n14451;
wire n14452;
wire n14453;
wire n14454;
wire n14455;
wire n14456;
wire n14457;
wire n14458;
wire n14459;
wire n14460;
wire n14461;
wire n14462;
wire n14463;
wire n14464;
wire n14465;
wire n14466;
wire n14467;
wire n14468;
wire n14469;
wire n14470;
wire n14471;
wire n14472;
wire n14473;
wire n14474;
wire n14475;
wire n14476;
wire n14477;
wire n14478;
wire n14479;
wire n14480;
wire n14481;
wire n14482;
wire n14483;
wire n14484;
wire n14485;
wire n14486;
wire n14487;
wire n14488;
wire n14489;
wire n14490;
wire n14491;
wire n14492;
wire n14493;
wire n14494;
wire n14495;
wire n14496;
wire n14497;
wire n14498;
wire n14499;
wire n14500;
wire n14501;
wire n14502;
wire n14503;
wire n14504;
wire n14505;
wire n14506;
wire n14507;
wire n14508;
wire n14509;
wire n14510;
wire n14511;
wire n14512;
wire n14513;
wire n14514;
wire n14515;
wire n14516;
wire n14517;
wire n14518;
wire n14519;
wire n14520;
wire n14521;
wire n14522;
wire n14523;
wire n14524;
wire n14525;
wire n14526;
wire n14527;
wire n14528;
wire n14529;
wire n14530;
wire n14531;
wire n14532;
wire n14533;
wire n14534;
wire n14535;
wire n14536;
wire n14537;
wire n14538;
wire n14539;
wire n14540;
wire n14541;
wire n14542;
wire n14543;
wire n14544;
wire n14545;
wire n14546;
wire n14547;
wire n14548;
wire n14549;
wire n14550;
wire n14551;
wire n14552;
wire n14553;
wire n14554;
wire n14555;
wire n14556;
wire n14557;
wire n14558;
wire n14559;
wire n14560;
wire n14561;
wire n14562;
wire n14563;
wire n14564;
wire n14565;
wire n14566;
wire n14567;
wire n14568;
wire n14569;
wire n14570;
wire n14571;
wire n14572;
wire n14573;
wire n14574;
wire n14575;
wire n14576;
wire n14577;
wire n14578;
wire n14579;
wire n14580;
wire n14581;
wire n14582;
wire n14583;
wire n14584;
wire n14585;
wire n14586;
wire n14587;
wire n14588;
wire n14589;
wire n14590;
wire n14591;
wire n14592;
wire n14593;
wire n14594;
wire n14595;
wire n14596;
wire n14597;
wire n14598;
wire n14599;
wire n14600;
wire n14601;
wire n14602;
wire n14603;
wire n14604;
wire n14605;
wire n14606;
wire n14607;
wire n14608;
wire n14609;
wire n14610;
wire n14611;
wire n14612;
wire n14613;
wire n14614;
wire n14615;
wire n14616;
wire n14617;
wire n14618;
wire n14619;
wire n14620;
wire n14621;
wire n14622;
wire n14623;
wire n14624;
wire n14625;
wire n14626;
wire n14627;
wire n14628;
wire n14629;
wire n14630;
wire n14631;
wire n14632;
wire n14633;
wire n14634;
wire n14635;
wire n14636;
wire n14637;
wire n14638;
wire n14639;
wire n14640;
wire n14641;
wire n14642;
wire n14643;
wire n14644;
wire n14645;
wire n14646;
wire n14647;
wire n14648;
wire n14649;
wire n14650;
wire n14651;
wire n14652;
wire n14653;
wire n14654;
wire n14655;
wire n14656;
wire n14657;
wire n14658;
wire n14659;
wire n14660;
wire n14661;
wire n14662;
wire n14663;
wire n14664;
wire n14665;
wire n14666;
wire n14667;
wire n14668;
wire n14669;
wire n14670;
wire n14671;
wire n14672;
wire n14673;
wire n14674;
wire n14675;
wire n14676;
wire n14677;
wire n14678;
wire n14679;
wire n14680;
wire n14681;
wire n14682;
wire n14683;
wire n14684;
wire n14685;
wire n14686;
wire n14687;
wire n14688;
wire n14689;
wire n14690;
wire n14691;
wire n14692;
wire n14693;
wire n14694;
wire n14695;
wire n14696;
wire n14697;
wire n14698;
wire n14699;
wire n14700;
wire n14701;
wire n14702;
wire n14703;
wire n14704;
wire n14705;
wire n14706;
wire n14707;
wire n14708;
wire n14709;
wire n14710;
wire n14711;
wire n14712;
wire n14713;
wire n14714;
wire n14715;
wire n14716;
wire n14717;
wire n14718;
wire n14719;
wire n14720;
wire n14721;
wire n14722;
wire n14723;
wire n14724;
wire n14725;
wire n14726;
wire n14727;
wire n14728;
wire n14729;
wire n14730;
wire n14731;
wire n14732;
wire n14733;
wire n14734;
wire n14735;
wire n14736;
wire n14737;
wire n14738;
wire n14739;
wire n14740;
wire n14741;
wire n14742;
wire n14743;
wire n14744;
wire n14745;
wire n14746;
wire n14747;
wire n14748;
wire n14749;
wire n14750;
wire n14751;
wire n14752;
wire n14753;
wire n14754;
wire n14755;
wire n14756;
wire n14757;
wire n14758;
wire n14759;
wire n14760;
wire n14761;
wire n14762;
wire n14763;
wire n14764;
wire n14765;
wire n14766;
wire n14767;
wire n14768;
wire n14769;
wire n14770;
wire n14771;
wire n14772;
wire n14773;
wire n14774;
wire n14775;
wire n14776;
wire n14777;
wire n14778;
wire n14779;
wire n14780;
wire n14781;
wire n14782;
wire n14783;
wire n14784;
wire n14785;
wire n14786;
wire n14787;
wire n14788;
wire n14789;
wire n14790;
wire n14791;
wire n14792;
wire n14793;
wire n14794;
wire n14795;
wire n14796;
wire n14797;
wire n14798;
wire n14799;
wire n14800;
wire n14801;
wire n14802;
wire n14803;
wire n14804;
wire n14805;
wire n14806;
wire n14807;
wire n14808;
wire n14809;
wire n14810;
wire n14811;
wire n14812;
wire n14813;
wire n14814;
wire n14815;
wire n14816;
wire n14817;
wire n14818;
wire n14819;
wire n14820;
wire n14821;
wire n14822;
wire n14823;
wire n14824;
wire n14825;
wire n14826;
wire n14827;
wire n14828;
wire n14829;
wire n14830;
wire n14831;
wire n14832;
wire n14833;
wire n14834;
wire n14835;
wire n14836;
wire n14837;
wire n14838;
wire n14839;
wire n14840;
wire n14841;
wire n14842;
wire n14843;
wire n14844;
wire n14845;
wire n14846;
wire n14847;
wire n14848;
wire n14849;
wire n14850;
wire n14851;
wire n14852;
wire n14853;
wire n14854;
wire n14855;
wire n14856;
wire n14857;
wire n14858;
wire n14859;
wire n14860;
wire n14861;
wire n14862;
wire n14863;
wire n14864;
wire n14865;
wire n14866;
wire n14867;
wire n14868;
wire n14869;
wire n14870;
wire n14871;
wire n14872;
wire n14873;
wire n14874;
wire n14875;
wire n14876;
wire n14877;
wire n14878;
wire n14879;
wire n14880;
wire n14881;
wire n14882;
wire n14883;
wire n14884;
wire n14885;
wire n14886;
wire n14887;
wire n14888;
wire n14889;
wire n14890;
wire n14891;
wire n14892;
wire n14893;
wire n14894;
wire n14895;
wire n14896;
wire n14897;
wire n14898;
wire n14899;
wire n14900;
wire n14901;
wire n14902;
wire n14903;
wire n14904;
wire n14905;
wire n14906;
wire n14907;
wire n14908;
wire n14909;
wire n14910;
wire n14911;
wire n14912;
wire n14913;
wire n14914;
wire n14915;
wire n14916;
wire n14917;
wire n14918;
wire n14919;
wire n14920;
wire n14921;
wire n14922;
wire n14923;
wire n14924;
wire n14925;
wire n14926;
wire n14927;
wire n14928;
wire n14929;
wire n14930;
wire n14931;
wire n14932;
wire n14933;
wire n14934;
wire n14935;
wire n14936;
wire n14937;
wire n14938;
wire n14939;
wire n14940;
wire n14941;
wire n14942;
wire n14943;
wire n14944;
wire n14945;
wire n14946;
wire n14947;
wire n14948;
wire n14949;
wire n14950;
wire n14951;
wire n14952;
wire n14953;
wire n14954;
wire n14955;
wire n14956;
wire n14957;
wire n14958;
wire n14959;
wire n14960;
wire n14961;
wire n14962;
wire n14963;
wire n14964;
wire n14965;
wire n14966;
wire n14967;
wire n14968;
wire n14969;
wire n14970;
wire n14971;
wire n14972;
wire n14973;
wire n14974;
wire n14975;
wire n14976;
wire n14977;
wire n14978;
wire n14979;
wire n14980;
wire n14981;
wire n14982;
wire n14983;
wire n14984;
wire n14985;
wire n14986;
wire n14987;
wire n14988;
wire n14989;
wire n14990;
wire n14991;
wire n14992;
wire n14993;
wire n14994;
wire n14995;
wire n14996;
wire n14997;
wire n14998;
wire n14999;
wire n15000;
wire n15001;
wire n15002;
wire n15003;
wire n15004;
wire n15005;
wire n15006;
wire n15007;
wire n15008;
wire n15009;
wire n15010;
wire n15011;
wire n15012;
wire n15013;
wire n15014;
wire n15015;
wire n15016;
wire n15017;
wire n15018;
wire n15019;
wire n15020;
wire n15021;
wire n15022;
wire n15023;
wire n15024;
wire n15025;
wire n15026;
wire n15027;
wire n15028;
wire n15029;
wire n15030;
wire n15031;
wire n15032;
wire n15033;
wire n15034;
wire n15035;
wire n15036;
wire n15037;
wire n15038;
wire n15039;
wire n15040;
wire n15041;
wire n15042;
wire n15043;
wire n15044;
wire n15045;
wire n15046;
wire n15047;
wire n15048;
wire n15049;
wire n15050;
wire n15051;
wire n15052;
wire n15053;
wire n15054;
wire n15055;
wire n15056;
wire n15057;
wire n15058;
wire n15059;
wire n15060;
wire n15061;
wire n15062;
wire n15063;
wire n15064;
wire n15065;
wire n15066;
wire n15067;
wire n15068;
wire n15069;
wire n15070;
wire n15071;
wire n15072;
wire n15073;
wire n15074;
wire n15075;
wire n15076;
wire n15077;
wire n15078;
wire n15079;
wire n15080;
wire n15081;
wire n15082;
wire n15083;
wire n15084;
wire n15085;
wire n15086;
wire n15087;
wire n15088;
wire n15089;
wire n15090;
wire n15091;
wire n15092;
wire n15093;
wire n15094;
wire n15095;
wire n15096;
wire n15097;
wire n15098;
wire n15099;
wire n15100;
wire n15101;
wire n15102;
wire n15103;
wire n15104;
wire n15105;
wire n15106;
wire n15107;
wire n15108;
wire n15109;
wire n15110;
wire n15111;
wire n15112;
wire n15113;
wire n15114;
wire n15115;
wire n15116;
wire n15117;
wire n15118;
wire n15119;
wire n15120;
wire n15121;
wire n15122;
wire n15123;
wire n15124;
wire n15125;
wire n15126;
wire n15127;
wire n15128;
wire n15129;
wire n15130;
wire n15131;
wire n15132;
wire n15133;
wire n15134;
wire n15135;
wire n15136;
wire n15137;
wire n15138;
wire n15139;
wire n15140;
wire n15141;
wire n15142;
wire n15143;
wire n15144;
wire n15145;
wire n15146;
wire n15147;
wire n15148;
wire n15149;
wire n15150;
wire n15151;
wire n15152;
wire n15153;
wire n15154;
wire n15155;
wire n15156;
wire n15157;
wire n15158;
wire n15159;
wire n15160;
wire n15161;
wire n15162;
wire n15163;
wire n15164;
wire n15165;
wire n15166;
wire n15167;
wire n15168;
wire n15169;
wire n15170;
wire n15171;
wire n15172;
wire n15173;
wire n15174;
wire n15175;
wire n15176;
wire n15177;
wire n15178;
wire n15179;
wire n15180;
wire n15181;
wire n15182;
wire n15183;
wire n15184;
wire n15185;
wire n15186;
wire n15187;
wire n15188;
wire n15189;
wire n15190;
wire n15191;
wire n15192;
wire n15193;
wire n15194;
wire n15195;
wire n15196;
wire n15197;
wire n15198;
wire n15199;
wire n15200;
wire n15201;
wire n15202;
wire n15203;
wire n15204;
wire n15205;
wire n15206;
wire n15207;
wire n15208;
wire n15209;
wire n15210;
wire n15211;
wire n15212;
wire n15213;
wire n15214;
wire n15215;
wire n15216;
wire n15217;
wire n15218;
wire n15219;
wire n15220;
wire n15221;
wire n15222;
wire n15223;
wire n15224;
wire n15225;
wire n15226;
wire n15227;
wire n15228;
wire n15229;
wire n15230;
wire n15231;
wire n15232;
wire n15233;
wire n15234;
wire n15235;
wire n15236;
wire n15237;
wire n15238;
wire n15239;
wire n15240;
wire n15241;
wire n15242;
wire n15243;
wire n15244;
wire n15245;
wire n15246;
wire n15247;
wire n15248;
wire n15249;
wire n15250;
wire n15251;
wire n15252;
wire n15253;
wire n15254;
wire n15255;
wire n15256;
wire n15257;
wire n15258;
wire n15259;
wire n15260;
wire n15261;
wire n15262;
wire n15263;
wire n15264;
wire n15265;
wire n15266;
wire n15267;
wire n15268;
wire n15269;
wire n15270;
wire n15271;
wire n15272;
wire n15273;
wire n15274;
wire n15275;
wire n15276;
wire n15277;
wire n15278;
wire n15279;
wire n15280;
wire n15281;
wire n15282;
wire n15283;
wire n15284;
wire n15285;
wire n15286;
wire n15287;
wire n15288;
wire n15289;
wire n15290;
wire n15291;
wire n15292;
wire n15293;
wire n15294;
wire n15295;
wire n15296;
wire n15297;
wire n15298;
wire n15299;
wire n15300;
wire n15301;
wire n15302;
wire n15303;
wire n15304;
wire n15305;
wire n15306;
wire n15307;
wire n15308;
wire n15309;
wire n15310;
wire n15311;
wire n15312;
wire n15313;
wire n15314;
wire n15315;
wire n15316;
wire n15317;
wire n15318;
wire n15319;
wire n15320;
wire n15321;
wire n15322;
wire n15323;
wire n15324;
wire n15325;
wire n15326;
wire n15327;
wire n15328;
wire n15329;
wire n15330;
wire n15331;
wire n15332;
wire n15333;
wire n15334;
wire n15335;
wire n15336;
wire n15337;
wire n15338;
wire n15339;
wire n15340;
wire n15341;
wire n15342;
wire n15343;
wire n15344;
wire n15345;
wire n15346;
wire n15347;
wire n15348;
wire n15349;
wire n15350;
wire n15351;
wire n15352;
wire n15353;
wire n15354;
wire n15355;
wire n15356;
wire n15357;
wire n15358;
wire n15359;
wire n15360;
wire n15361;
wire n15362;
wire n15363;
wire n15364;
wire n15365;
wire n15366;
wire n15367;
wire n15368;
wire n15369;
wire n15370;
wire n15371;
wire n15372;
wire n15373;
wire n15374;
wire n15375;
wire n15376;
wire n15377;
wire n15378;
wire n15379;
wire n15380;
wire n15381;
wire n15382;
wire n15383;
wire n15384;
wire n15385;
wire n15386;
wire n15387;
wire n15388;
wire n15389;
wire n15390;
wire n15391;
wire n15392;
wire n15393;
wire n15394;
wire n15395;
wire n15396;
wire n15397;
wire n15398;
wire n15399;
wire n15400;
wire n15401;
wire n15402;
wire n15403;
wire n15404;
wire n15405;
wire n15406;
wire n15407;
wire n15408;
wire n15409;
wire n15410;
wire n15411;
wire n15412;
wire n15413;
wire n15414;
wire n15415;
wire n15416;
wire n15417;
wire n15418;
wire n15419;
wire n15420;
wire n15421;
wire n15422;
wire n15423;
wire n15424;
wire n15425;
wire n15426;
wire n15427;
wire n15428;
wire n15429;
wire n15430;
wire n15431;
wire n15432;
wire n15433;
wire n15434;
wire n15435;
wire n15436;
wire n15437;
wire n15438;
wire n15439;
wire n15440;
wire n15441;
wire n15442;
wire n15443;
wire n15444;
wire n15445;
wire n15446;
wire n15447;
wire n15448;
wire n15449;
wire n15450;
wire n15451;
wire n15452;
wire n15453;
wire n15454;
wire n15455;
wire n15456;
wire n15457;
wire n15458;
wire n15459;
wire n15460;
wire n15461;
wire n15462;
wire n15463;
wire n15464;
wire n15465;
wire n15466;
wire n15467;
wire n15468;
wire n15469;
wire n15470;
wire n15471;
wire n15472;
wire n15473;
wire n15474;
wire n15475;
wire n15476;
wire n15477;
wire n15478;
wire n15479;
wire n15480;
wire n15481;
wire n15482;
wire n15483;
wire n15484;
wire n15485;
wire n15486;
wire n15487;
wire n15488;
wire n15489;
wire n15490;
wire n15491;
wire n15492;
wire n15493;
wire n15494;
wire n15495;
wire n15496;
wire n15497;
wire n15498;
wire n15499;
wire n15500;
wire n15501;
wire n15502;
wire n15503;
wire n15504;
wire n15505;
wire n15506;
wire n15507;
wire n15508;
wire n15509;
wire n15510;
wire n15511;
wire n15512;
wire n15513;
wire n15514;
wire n15515;
wire n15516;
wire n15517;
wire n15518;
wire n15519;
wire n15520;
wire n15521;
wire n15522;
wire n15523;
wire _i_CLEFIA128_keyL_0;
wire _i_CLEFIA128_keyL_1;
wire _i_CLEFIA128_keyL_2;
wire _i_CLEFIA128_keyL_3;
wire _i_CLEFIA128_keyL_4;
wire _i_CLEFIA128_keyL_5;
wire _i_CLEFIA128_keyL_6;
wire _i_CLEFIA128_keyL_7;
wire _i_CLEFIA128_keyL_8;
wire _i_CLEFIA128_keyL_9;
wire _i_CLEFIA128_keyL_10;
wire _i_CLEFIA128_keyL_11;
wire _i_CLEFIA128_keyL_12;
wire _i_CLEFIA128_keyL_13;
wire _i_CLEFIA128_keyL_14;
wire _i_CLEFIA128_keyL_15;
wire _i_CLEFIA128_keyL_16;
wire _i_CLEFIA128_keyL_17;
wire _i_CLEFIA128_keyL_18;
wire _i_CLEFIA128_keyL_19;
wire _i_CLEFIA128_keyL_20;
wire _i_CLEFIA128_keyL_21;
wire _i_CLEFIA128_keyL_22;
wire _i_CLEFIA128_keyL_23;
wire _i_CLEFIA128_keyL_24;
wire _i_CLEFIA128_keyL_25;
wire _i_CLEFIA128_keyL_26;
wire _i_CLEFIA128_keyL_27;
wire _i_CLEFIA128_keyL_28;
wire _i_CLEFIA128_keyL_29;
wire _i_CLEFIA128_keyL_30;
wire _i_CLEFIA128_keyL_31;
wire _i_CLEFIA128_keyL_32;
wire _i_CLEFIA128_keyL_33;
wire _i_CLEFIA128_keyL_34;
wire _i_CLEFIA128_keyL_35;
wire _i_CLEFIA128_keyL_36;
wire _i_CLEFIA128_keyL_37;
wire _i_CLEFIA128_keyL_38;
wire _i_CLEFIA128_keyL_39;
wire _i_CLEFIA128_keyL_40;
wire _i_CLEFIA128_keyL_41;
wire _i_CLEFIA128_keyL_42;
wire _i_CLEFIA128_keyL_43;
wire _i_CLEFIA128_keyL_44;
wire _i_CLEFIA128_keyL_45;
wire _i_CLEFIA128_keyL_46;
wire _i_CLEFIA128_keyL_47;
wire _i_CLEFIA128_keyL_48;
wire _i_CLEFIA128_keyL_49;
wire _i_CLEFIA128_keyL_50;
wire _i_CLEFIA128_keyL_51;
wire _i_CLEFIA128_keyL_52;
wire _i_CLEFIA128_keyL_53;
wire _i_CLEFIA128_keyL_54;
wire _i_CLEFIA128_keyL_55;
wire _i_CLEFIA128_keyL_56;
wire _i_CLEFIA128_keyL_57;
wire _i_CLEFIA128_keyL_58;
wire _i_CLEFIA128_keyL_59;
wire _i_CLEFIA128_keyL_60;
wire _i_CLEFIA128_keyL_61;
wire _i_CLEFIA128_keyL_62;
wire _i_CLEFIA128_keyL_63;
wire _i_CLEFIA128_keyL_64;
wire _i_CLEFIA128_keyL_65;
wire _i_CLEFIA128_keyL_66;
wire _i_CLEFIA128_keyL_67;
wire _i_CLEFIA128_keyL_68;
wire _i_CLEFIA128_keyL_69;
wire _i_CLEFIA128_keyL_70;
wire _i_CLEFIA128_keyL_71;
wire _i_CLEFIA128_keyL_72;
wire _i_CLEFIA128_keyL_73;
wire _i_CLEFIA128_keyL_74;
wire _i_CLEFIA128_keyL_75;
wire _i_CLEFIA128_keyL_76;
wire _i_CLEFIA128_keyL_77;
wire _i_CLEFIA128_keyL_78;
wire _i_CLEFIA128_keyL_79;
wire _i_CLEFIA128_keyL_80;
wire _i_CLEFIA128_keyL_81;
wire _i_CLEFIA128_keyL_82;
wire _i_CLEFIA128_keyL_83;
wire _i_CLEFIA128_keyL_84;
wire _i_CLEFIA128_keyL_85;
wire _i_CLEFIA128_keyL_86;
wire _i_CLEFIA128_keyL_87;
wire _i_CLEFIA128_keyL_88;
wire _i_CLEFIA128_keyL_89;
wire _i_CLEFIA128_keyL_90;
wire _i_CLEFIA128_keyL_91;
wire _i_CLEFIA128_keyL_92;
wire _i_CLEFIA128_keyL_93;
wire _i_CLEFIA128_keyL_94;
wire _i_CLEFIA128_keyL_95;
wire _i_CLEFIA128_keyL_96;
wire _i_CLEFIA128_keyL_97;
wire _i_CLEFIA128_keyL_98;
wire _i_CLEFIA128_keyL_99;
wire _i_CLEFIA128_keyL_100;
wire _i_CLEFIA128_keyL_101;
wire _i_CLEFIA128_keyL_102;
wire _i_CLEFIA128_keyL_103;
wire _i_CLEFIA128_keyL_104;
wire _i_CLEFIA128_keyL_105;
wire _i_CLEFIA128_keyL_106;
wire _i_CLEFIA128_keyL_107;
wire _i_CLEFIA128_keyL_108;
wire _i_CLEFIA128_keyL_109;
wire _i_CLEFIA128_keyL_110;
wire _i_CLEFIA128_keyL_111;
wire _i_CLEFIA128_keyL_112;
wire _i_CLEFIA128_keyL_113;
wire _i_CLEFIA128_keyL_114;
wire _i_CLEFIA128_keyL_115;
wire _i_CLEFIA128_keyL_116;
wire _i_CLEFIA128_keyL_117;
wire _i_CLEFIA128_keyL_118;
wire _i_CLEFIA128_keyL_119;
wire _i_CLEFIA128_keyL_120;
wire _i_CLEFIA128_keyL_121;
wire _i_CLEFIA128_keyL_122;
wire _i_CLEFIA128_keyL_123;
wire _i_CLEFIA128_keyL_124;
wire _i_CLEFIA128_keyL_125;
wire _i_CLEFIA128_keyL_126;
wire _i_CLEFIA128_keyL_127;
wire _i_CLEFIA128_keyK_0;
wire _i_CLEFIA128_keyK_1;
wire _i_CLEFIA128_keyK_2;
wire _i_CLEFIA128_keyK_3;
wire _i_CLEFIA128_keyK_4;
wire _i_CLEFIA128_keyK_5;
wire _i_CLEFIA128_keyK_6;
wire _i_CLEFIA128_keyK_7;
wire _i_CLEFIA128_keyK_8;
wire _i_CLEFIA128_keyK_9;
wire _i_CLEFIA128_keyK_10;
wire _i_CLEFIA128_keyK_11;
wire _i_CLEFIA128_keyK_12;
wire _i_CLEFIA128_keyK_13;
wire _i_CLEFIA128_keyK_14;
wire _i_CLEFIA128_keyK_15;
wire _i_CLEFIA128_keyK_16;
wire _i_CLEFIA128_keyK_17;
wire _i_CLEFIA128_keyK_18;
wire _i_CLEFIA128_keyK_19;
wire _i_CLEFIA128_keyK_20;
wire _i_CLEFIA128_keyK_21;
wire _i_CLEFIA128_keyK_22;
wire _i_CLEFIA128_keyK_23;
wire _i_CLEFIA128_keyK_24;
wire _i_CLEFIA128_keyK_25;
wire _i_CLEFIA128_keyK_26;
wire _i_CLEFIA128_keyK_27;
wire _i_CLEFIA128_keyK_28;
wire _i_CLEFIA128_keyK_29;
wire _i_CLEFIA128_keyK_30;
wire _i_CLEFIA128_keyK_31;
wire _i_CLEFIA128_keyK_32;
wire _i_CLEFIA128_keyK_33;
wire _i_CLEFIA128_keyK_34;
wire _i_CLEFIA128_keyK_35;
wire _i_CLEFIA128_keyK_36;
wire _i_CLEFIA128_keyK_37;
wire _i_CLEFIA128_keyK_38;
wire _i_CLEFIA128_keyK_39;
wire _i_CLEFIA128_keyK_40;
wire _i_CLEFIA128_keyK_41;
wire _i_CLEFIA128_keyK_42;
wire _i_CLEFIA128_keyK_43;
wire _i_CLEFIA128_keyK_44;
wire _i_CLEFIA128_keyK_45;
wire _i_CLEFIA128_keyK_46;
wire _i_CLEFIA128_keyK_47;
wire _i_CLEFIA128_keyK_48;
wire _i_CLEFIA128_keyK_49;
wire _i_CLEFIA128_keyK_50;
wire _i_CLEFIA128_keyK_51;
wire _i_CLEFIA128_keyK_52;
wire _i_CLEFIA128_keyK_53;
wire _i_CLEFIA128_keyK_54;
wire _i_CLEFIA128_keyK_55;
wire _i_CLEFIA128_keyK_56;
wire _i_CLEFIA128_keyK_57;
wire _i_CLEFIA128_keyK_58;
wire _i_CLEFIA128_keyK_59;
wire _i_CLEFIA128_keyK_60;
wire _i_CLEFIA128_keyK_61;
wire _i_CLEFIA128_keyK_62;
wire _i_CLEFIA128_keyK_63;
wire _i_CLEFIA128_keyK_64;
wire _i_CLEFIA128_keyK_65;
wire _i_CLEFIA128_keyK_66;
wire _i_CLEFIA128_keyK_67;
wire _i_CLEFIA128_keyK_68;
wire _i_CLEFIA128_keyK_69;
wire _i_CLEFIA128_keyK_70;
wire _i_CLEFIA128_keyK_71;
wire _i_CLEFIA128_keyK_72;
wire _i_CLEFIA128_keyK_73;
wire _i_CLEFIA128_keyK_74;
wire _i_CLEFIA128_keyK_75;
wire _i_CLEFIA128_keyK_76;
wire _i_CLEFIA128_keyK_77;
wire _i_CLEFIA128_keyK_78;
wire _i_CLEFIA128_keyK_79;
wire _i_CLEFIA128_keyK_80;
wire _i_CLEFIA128_keyK_81;
wire _i_CLEFIA128_keyK_82;
wire _i_CLEFIA128_keyK_83;
wire _i_CLEFIA128_keyK_84;
wire _i_CLEFIA128_keyK_85;
wire _i_CLEFIA128_keyK_86;
wire _i_CLEFIA128_keyK_87;
wire _i_CLEFIA128_keyK_88;
wire _i_CLEFIA128_keyK_89;
wire _i_CLEFIA128_keyK_90;
wire _i_CLEFIA128_keyK_91;
wire _i_CLEFIA128_keyK_92;
wire _i_CLEFIA128_keyK_93;
wire _i_CLEFIA128_keyK_94;
wire _i_CLEFIA128_keyK_95;
wire _i_CLEFIA128_keyK_96;
wire _i_CLEFIA128_keyK_97;
wire _i_CLEFIA128_keyK_98;
wire _i_CLEFIA128_keyK_99;
wire _i_CLEFIA128_keyK_100;
wire _i_CLEFIA128_keyK_101;
wire _i_CLEFIA128_keyK_102;
wire _i_CLEFIA128_keyK_103;
wire _i_CLEFIA128_keyK_104;
wire _i_CLEFIA128_keyK_105;
wire _i_CLEFIA128_keyK_106;
wire _i_CLEFIA128_keyK_107;
wire _i_CLEFIA128_keyK_108;
wire _i_CLEFIA128_keyK_109;
wire _i_CLEFIA128_keyK_110;
wire _i_CLEFIA128_keyK_111;
wire _i_CLEFIA128_keyK_112;
wire _i_CLEFIA128_keyK_113;
wire _i_CLEFIA128_keyK_114;
wire _i_CLEFIA128_keyK_115;
wire _i_CLEFIA128_keyK_116;
wire _i_CLEFIA128_keyK_117;
wire _i_CLEFIA128_keyK_118;
wire _i_CLEFIA128_keyK_119;
wire _i_CLEFIA128_keyK_120;
wire _i_CLEFIA128_keyK_121;
wire _i_CLEFIA128_keyK_122;
wire _i_CLEFIA128_keyK_123;
wire _i_CLEFIA128_keyK_124;
wire _i_CLEFIA128_keyK_125;
wire _i_CLEFIA128_keyK_126;
wire _i_CLEFIA128_keyK_127;
wire _i_CLEFIA128_CON_T_xi_9;
wire _i_CLEFIA128_CON_T_xi_10;
wire _i_CLEFIA128_CON_T_xi_11;
wire _i_CLEFIA128_CON_T_xi_12;
wire _i_CLEFIA128_CON_T_xi_13;
wire _i_CLEFIA128_CON_T_xi_14;
wire _i_CLEFIA128_CON_T_x_0;
wire _i_CLEFIA128_CON_T_x_1;
wire _i_CLEFIA128_CON_T_x_2;
wire _i_CLEFIA128_CON_T_x_3;
wire _i_CLEFIA128_CON_T_x_4;
wire _i_CLEFIA128_CON_T_x_5;
wire _i_CLEFIA128_CON_T_x_6;
wire _i_CLEFIA128_CON_T_x_7;
wire _i_CLEFIA128_CON_T_x_8;
wire _i_CLEFIA128_CON_T_x_9;
wire _i_CLEFIA128_CON_T_x_10;
wire _i_CLEFIA128_CON_T_x_11;
wire _i_CLEFIA128_CON_T_x_12;
wire _i_CLEFIA128_CON_T_x_13;
wire _i_CLEFIA128_CON_T_x_14;
wire _i_CLEFIA128_CON_T_x_15;
wire _i_CLEFIA128_rndcnt_reg_0;
wire _i_CLEFIA128_rndcnt_reg_1;
wire _i_CLEFIA128_rndcnt_reg_2;
wire _i_CLEFIA128_rndcnt_reg_3;
wire _i_CLEFIA128_rndcnt_reg_4;
wire _i_CLEFIA128_state_reg_0;
wire _i_CLEFIA128_state_reg_1;
//Start cells  
  QDFFHHD _i_CLEFIA128_BSY_reg_reg  ( .D(n6503), .CK(CLK), .Q(BSY) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_0  ( .D(n6502), .CK(CLK), .Q(_i_CLEFIA128_keyK _0) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_29  ( .D(n6501), .CK(CLK), .Q(_i_CLEFIA128_keyK _29) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_30  ( .D(n6500), .CK(CLK), .Q(_i_CLEFIA128_keyK _30) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_31  ( .D(n6499), .CK(CLK), .Q(_i_CLEFIA128_keyK _31) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_32  ( .D(n6498), .CK(CLK), .Q(_i_CLEFIA128_keyK _32) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_33  ( .D(n6497), .CK(CLK), .Q(_i_CLEFIA128_keyK _33) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_34  ( .D(n6496), .CK(CLK), .Q(_i_CLEFIA128_keyK _34) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_35  ( .D(n6495), .CK(CLK), .Q(_i_CLEFIA128_keyK _35) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_36  ( .D(n6494), .CK(CLK), .Q(_i_CLEFIA128_keyK _36) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_37  ( .D(n6493), .CK(CLK), .Q(_i_CLEFIA128_keyK _37) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_38  ( .D(n6492), .CK(CLK), .Q(_i_CLEFIA128_keyK _38) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_39  ( .D(n6491), .CK(CLK), .Q(_i_CLEFIA128_keyK _39) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_40  ( .D(n6490), .CK(CLK), .Q(_i_CLEFIA128_keyK _40) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_41  ( .D(n6489), .CK(CLK), .Q(_i_CLEFIA128_keyK _41) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_42  ( .D(n6488), .CK(CLK), .Q(_i_CLEFIA128_keyK _42) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_43  ( .D(n6487), .CK(CLK), .Q(_i_CLEFIA128_keyK _43) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_44  ( .D(n6486), .CK(CLK), .Q(_i_CLEFIA128_keyK _44) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_45  ( .D(n6485), .CK(CLK), .Q(_i_CLEFIA128_keyK _45) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_46  ( .D(n6484), .CK(CLK), .Q(_i_CLEFIA128_keyK _46) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_47  ( .D(n6483), .CK(CLK), .Q(_i_CLEFIA128_keyK _47) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_48  ( .D(n6482), .CK(CLK), .Q(_i_CLEFIA128_keyK _48) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_49  ( .D(n6481), .CK(CLK), .Q(_i_CLEFIA128_keyK _49) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_50  ( .D(n6480), .CK(CLK), .Q(_i_CLEFIA128_keyK _50) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_51  ( .D(n6479), .CK(CLK), .Q(_i_CLEFIA128_keyK _51) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_52  ( .D(n6478), .CK(CLK), .Q(_i_CLEFIA128_keyK _52) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_53  ( .D(n6477), .CK(CLK), .Q(_i_CLEFIA128_keyK _53) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_54  ( .D(n6476), .CK(CLK), .Q(_i_CLEFIA128_keyK _54) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_55  ( .D(n6475), .CK(CLK), .Q(_i_CLEFIA128_keyK _55) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_56  ( .D(n6474), .CK(CLK), .Q(_i_CLEFIA128_keyK _56) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_57  ( .D(n6473), .CK(CLK), .Q(_i_CLEFIA128_keyK _57) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_58  ( .D(n6472), .CK(CLK), .Q(_i_CLEFIA128_keyK _58) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_59  ( .D(n6471), .CK(CLK), .Q(_i_CLEFIA128_keyK _59) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_60  ( .D(n6470), .CK(CLK), .Q(_i_CLEFIA128_keyK _60) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_61  ( .D(n6469), .CK(CLK), .Q(_i_CLEFIA128_keyK _61) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_62  ( .D(n6468), .CK(CLK), .Q(_i_CLEFIA128_keyK _62) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_63  ( .D(n6467), .CK(CLK), .Q(_i_CLEFIA128_keyK _63) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_64  ( .D(n6466), .CK(CLK), .Q(_i_CLEFIA128_keyK _64) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_65  ( .D(n6465), .CK(CLK), .Q(_i_CLEFIA128_keyK _65) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_66  ( .D(n6464), .CK(CLK), .Q(_i_CLEFIA128_keyK _66) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_67  ( .D(n6463), .CK(CLK), .Q(_i_CLEFIA128_keyK _67) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_68  ( .D(n6462), .CK(CLK), .Q(_i_CLEFIA128_keyK _68) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_69  ( .D(n6461), .CK(CLK), .Q(_i_CLEFIA128_keyK _69) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_70  ( .D(n6460), .CK(CLK), .Q(_i_CLEFIA128_keyK _70) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_71  ( .D(n6459), .CK(CLK), .Q(_i_CLEFIA128_keyK _71) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_72  ( .D(n6458), .CK(CLK), .Q(_i_CLEFIA128_keyK _72) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_73  ( .D(n6457), .CK(CLK), .Q(_i_CLEFIA128_keyK _73) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_74  ( .D(n6456), .CK(CLK), .Q(_i_CLEFIA128_keyK _74) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_75  ( .D(n6455), .CK(CLK), .Q(_i_CLEFIA128_keyK _75) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_76  ( .D(n6454), .CK(CLK), .Q(_i_CLEFIA128_keyK _76) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_77  ( .D(n6453), .CK(CLK), .Q(_i_CLEFIA128_keyK _77) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_78  ( .D(n6452), .CK(CLK), .Q(_i_CLEFIA128_keyK _78) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_79  ( .D(n6451), .CK(CLK), .Q(_i_CLEFIA128_keyK _79) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_80  ( .D(n6450), .CK(CLK), .Q(_i_CLEFIA128_keyK _80) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_81  ( .D(n6449), .CK(CLK), .Q(_i_CLEFIA128_keyK _81) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_82  ( .D(n6448), .CK(CLK), .Q(_i_CLEFIA128_keyK _82) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_83  ( .D(n6447), .CK(CLK), .Q(_i_CLEFIA128_keyK _83) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_84  ( .D(n6446), .CK(CLK), .Q(_i_CLEFIA128_keyK _84) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_85  ( .D(n6445), .CK(CLK), .Q(_i_CLEFIA128_keyK _85) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_86  ( .D(n6444), .CK(CLK), .Q(_i_CLEFIA128_keyK _86) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_87  ( .D(n6443), .CK(CLK), .Q(_i_CLEFIA128_keyK _87) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_88  ( .D(n6442), .CK(CLK), .Q(_i_CLEFIA128_keyK _88) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_89  ( .D(n6441), .CK(CLK), .Q(_i_CLEFIA128_keyK _89) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_90  ( .D(n6440), .CK(CLK), .Q(_i_CLEFIA128_keyK _90) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_91  ( .D(n6439), .CK(CLK), .Q(_i_CLEFIA128_keyK _91) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_92  ( .D(n6438), .CK(CLK), .Q(_i_CLEFIA128_keyK _92) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_93  ( .D(n6437), .CK(CLK), .Q(_i_CLEFIA128_keyK _93) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_94  ( .D(n6436), .CK(CLK), .Q(_i_CLEFIA128_keyK _94) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_95  ( .D(n6435), .CK(CLK), .Q(_i_CLEFIA128_keyK _95) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_96  ( .D(n6434), .CK(CLK), .Q(_i_CLEFIA128_keyK _96) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_97  ( .D(n6433), .CK(CLK), .Q(_i_CLEFIA128_keyK _97) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_98  ( .D(n6432), .CK(CLK), .Q(_i_CLEFIA128_keyK _98) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_99  ( .D(n6431), .CK(CLK), .Q(_i_CLEFIA128_keyK _99) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_100  ( .D(n6430), .CK(CLK), .Q(_i_CLEFIA128_keyK _100) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_101  ( .D(n6429), .CK(CLK), .Q(_i_CLEFIA128_keyK _101) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_102  ( .D(n6428), .CK(CLK), .Q(_i_CLEFIA128_keyK _102) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_103  ( .D(n6427), .CK(CLK), .Q(_i_CLEFIA128_keyK _103) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_104  ( .D(n6426), .CK(CLK), .Q(_i_CLEFIA128_keyK _104) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_105  ( .D(n6425), .CK(CLK), .Q(_i_CLEFIA128_keyK _105) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_106  ( .D(n6424), .CK(CLK), .Q(_i_CLEFIA128_keyK _106) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_107  ( .D(n6423), .CK(CLK), .Q(_i_CLEFIA128_keyK _107) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_108  ( .D(n6422), .CK(CLK), .Q(_i_CLEFIA128_keyK _108) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_109  ( .D(n6421), .CK(CLK), .Q(_i_CLEFIA128_keyK _109) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_110  ( .D(n6420), .CK(CLK), .Q(_i_CLEFIA128_keyK _110) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_111  ( .D(n6419), .CK(CLK), .Q(_i_CLEFIA128_keyK _111) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_112  ( .D(n6418), .CK(CLK), .Q(_i_CLEFIA128_keyK _112) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_113  ( .D(n6417), .CK(CLK), .Q(_i_CLEFIA128_keyK _113) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_114  ( .D(n6416), .CK(CLK), .Q(_i_CLEFIA128_keyK _114) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_115  ( .D(n6415), .CK(CLK), .Q(_i_CLEFIA128_keyK _115) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_116  ( .D(n6414), .CK(CLK), .Q(_i_CLEFIA128_keyK _116) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_117  ( .D(n6413), .CK(CLK), .Q(_i_CLEFIA128_keyK _117) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_118  ( .D(n6412), .CK(CLK), .Q(_i_CLEFIA128_keyK _118) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_119  ( .D(n6411), .CK(CLK), .Q(_i_CLEFIA128_keyK _119) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_120  ( .D(n6410), .CK(CLK), .Q(_i_CLEFIA128_keyK _120) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_121  ( .D(n6409), .CK(CLK), .Q(_i_CLEFIA128_keyK _121) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_122  ( .D(n6408), .CK(CLK), .Q(_i_CLEFIA128_keyK _122) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_123  ( .D(n6407), .CK(CLK), .Q(_i_CLEFIA128_keyK _123) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_124  ( .D(n6406), .CK(CLK), .Q(_i_CLEFIA128_keyK _124) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_125  ( .D(n6405), .CK(CLK), .Q(_i_CLEFIA128_keyK _125) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_126  ( .D(n6404), .CK(CLK), .Q(_i_CLEFIA128_keyK _126) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_127  ( .D(n6403), .CK(CLK), .Q(_i_CLEFIA128_keyK _127) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_1  ( .D(n6402), .CK(CLK), .Q(_i_CLEFIA128_keyK _1) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_2  ( .D(n6401), .CK(CLK), .Q(_i_CLEFIA128_keyK _2) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_3  ( .D(n6400), .CK(CLK), .Q(_i_CLEFIA128_keyK _3) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_4  ( .D(n6399), .CK(CLK), .Q(_i_CLEFIA128_keyK _4) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_5  ( .D(n6398), .CK(CLK), .Q(_i_CLEFIA128_keyK _5) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_6  ( .D(n6397), .CK(CLK), .Q(_i_CLEFIA128_keyK _6) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_7  ( .D(n6396), .CK(CLK), .Q(_i_CLEFIA128_keyK _7) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_8  ( .D(n6395), .CK(CLK), .Q(_i_CLEFIA128_keyK _8) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_9  ( .D(n6394), .CK(CLK), .Q(_i_CLEFIA128_keyK _9) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_10  ( .D(n6393), .CK(CLK), .Q(_i_CLEFIA128_keyK _10) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_11  ( .D(n6392), .CK(CLK), .Q(_i_CLEFIA128_keyK _11) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_12  ( .D(n6391), .CK(CLK), .Q(_i_CLEFIA128_keyK _12) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_13  ( .D(n6390), .CK(CLK), .Q(_i_CLEFIA128_keyK _13) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_14  ( .D(n6389), .CK(CLK), .Q(_i_CLEFIA128_keyK _14) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_15  ( .D(n6388), .CK(CLK), .Q(_i_CLEFIA128_keyK _15) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_16  ( .D(n6387), .CK(CLK), .Q(_i_CLEFIA128_keyK _16) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_17  ( .D(n6386), .CK(CLK), .Q(_i_CLEFIA128_keyK _17) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_18  ( .D(n6385), .CK(CLK), .Q(_i_CLEFIA128_keyK _18) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_19  ( .D(n6384), .CK(CLK), .Q(_i_CLEFIA128_keyK _19) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_20  ( .D(n6383), .CK(CLK), .Q(_i_CLEFIA128_keyK _20) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_21  ( .D(n6382), .CK(CLK), .Q(_i_CLEFIA128_keyK _21) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_22  ( .D(n6381), .CK(CLK), .Q(_i_CLEFIA128_keyK _22) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_23  ( .D(n6380), .CK(CLK), .Q(_i_CLEFIA128_keyK _23) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_24  ( .D(n6379), .CK(CLK), .Q(_i_CLEFIA128_keyK _24) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_25  ( .D(n6378), .CK(CLK), .Q(_i_CLEFIA128_keyK _25) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_26  ( .D(n6377), .CK(CLK), .Q(_i_CLEFIA128_keyK _26) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_27  ( .D(n6376), .CK(CLK), .Q(_i_CLEFIA128_keyK _27) );
  QDFFHHD _i_CLEFIA128_keyK_reg_reg_28  ( .D(n6375), .CK(CLK), .Q(_i_CLEFIA128_keyK _28) );
  QDFFHHD _i_CLEFIA128_state_reg_reg_0  ( .D(n6368), .CK(CLK), .Q(_i_CLEFIA128_state_reg _0) );
  QDFFHHD _i_CLEFIA128_state_reg_reg_1  ( .D(n6367), .CK(CLK), .Q(_i_CLEFIA128_state_reg _1) );
  QDFFHHD _i_CLEFIA128_rndcnt_reg_reg_2  ( .D(n6371), .CK(CLK), .Q(_i_CLEFIA128_rndcnt_reg _2) );
  QDFFHHD _i_CLEFIA128_rndcnt_reg_reg_3  ( .D(n6372), .CK(CLK), .Q(_i_CLEFIA128_rndcnt_reg _3) );
  QDFFHHD _i_CLEFIA128_rndcnt_reg_reg_4  ( .D(n6373), .CK(CLK), .Q(_i_CLEFIA128_rndcnt_reg _4) );
  QDFFHHD _i_CLEFIA128_rndcnt_reg_reg_0  ( .D(n6374), .CK(CLK), .Q(_i_CLEFIA128_rndcnt_reg _0) );
  QDFFHHD _i_CLEFIA128_CON_T_reg_reg_14  ( .D(n6351), .CK(CLK), .Q(_i_CLEFIA128_CON_T_xi _13) );
  QDFFHHD _i_CLEFIA128_CON_T_reg_reg_13  ( .D(n6352), .CK(CLK), .Q(_i_CLEFIA128_CON_T_x _14) );
  QDFFHHD _i_CLEFIA128_CON_T_reg_reg_12  ( .D(n6353), .CK(CLK), .Q(_i_CLEFIA128_CON_T_xi _11) );
  QDFFHHD _i_CLEFIA128_CON_T_reg_reg_11  ( .D(n6354), .CK(CLK), .Q(_i_CLEFIA128_CON_T_x _12) );
  QDFFHHD _i_CLEFIA128_CON_T_reg_reg_10  ( .D(n6355), .CK(CLK), .Q(_i_CLEFIA128_CON_T_xi _9) );
  QDFFHHD _i_CLEFIA128_CON_T_reg_reg_9  ( .D(n6356), .CK(CLK), .Q(_i_CLEFIA128_CON_T_x _10) );
  QDFFHHD _i_CLEFIA128_CON_T_reg_reg_8  ( .D(n6357), .CK(CLK), .Q(_i_CLEFIA128_CON_T_x _9) );
  QDFFHHD _i_CLEFIA128_CON_T_reg_reg_7  ( .D(n6358), .CK(CLK), .Q(_i_CLEFIA128_CON_T_x _8) );
  QDFFHHD _i_CLEFIA128_CON_T_reg_reg_6  ( .D(n6359), .CK(CLK), .Q(_i_CLEFIA128_CON_T_x _7) );
  QDFFHHD _i_CLEFIA128_CON_T_reg_reg_5  ( .D(n6360), .CK(CLK), .Q(_i_CLEFIA128_CON_T_x _6) );
  QDFFHHD _i_CLEFIA128_CON_T_reg_reg_4  ( .D(n6361), .CK(CLK), .Q(_i_CLEFIA128_CON_T_reg_4 ) );
  QDFFHHD _i_CLEFIA128_CON_T_reg_reg_3  ( .D(n6362), .CK(CLK), .Q(_i_CLEFIA128_CON_T_xi_2 ) );
  QDFFHHD _i_CLEFIA128_CON_T_reg_reg_2  ( .D(n6363), .CK(CLK), .Q(_i_CLEFIA128_CON_T_x _3) );
  QDFFHHD _i_CLEFIA128_CON_T_reg_reg_1  ( .D(n6364), .CK(CLK), .Q(_i_CLEFIA128_CON_T_x _2) );
  QDFFHHD _i_CLEFIA128_CON_T_reg_reg_0  ( .D(n6365), .CK(CLK), .Q(_i_CLEFIA128_CON_T_x _1) );
  QDFFHHD _i_CLEFIA128_CON_T_reg_reg_15  ( .D(n6366), .CK(CLK), .Q(_i_CLEFIA128_CON_T_x _0) );
  QDFFHHD _i_CLEFIA128_data1_reg_reg_0  ( .D(n6095), .CK(CLK), .Q(DOUT_64));
  QDFFHHD _i_CLEFIA128_data0_reg_reg_0  ( .D(n6190), .CK(CLK), .Q(DOUT_96));
  QDFFHHD _i_CLEFIA128_data2_reg_reg_26  ( .D(n6184), .CK(CLK), .Q(DOUT_58));
  QDFFHHD _i_CLEFIA128_data2_reg_reg_31  ( .D(n6189), .CK(CLK), .Q(DOUT_63));
  QDFFHHD _i_CLEFIA128_data2_reg_reg_30  ( .D(n6188), .CK(CLK), .Q(DOUT_62));
  QDFFHHD _i_CLEFIA128_data2_reg_reg_29  ( .D(n6187), .CK(CLK), .Q(DOUT_61));
  QDFFHHD _i_CLEFIA128_data2_reg_reg_24  ( .D(n6182), .CK(CLK), .Q(DOUT_56));
  QDFFHHD _i_CLEFIA128_data2_reg_reg_27  ( .D(n6185), .CK(CLK), .Q(DOUT_59));
  QDFFHHD _i_CLEFIA128_data2_reg_reg_28  ( .D(n6186), .CK(CLK), .Q(DOUT_60));
  QDFFHHD _i_CLEFIA128_data0_reg_reg_26  ( .D(n6216), .CK(CLK), .Q(DOUT_122));
  QDFFHHD _i_CLEFIA128_data2_reg_reg_12  ( .D(n6170), .CK(CLK), .Q(DOUT_44));
  QDFFHHD _i_CLEFIA128_data2_reg_reg_23  ( .D(n6181), .CK(CLK), .Q(DOUT_55));
  QDFFHHD _i_CLEFIA128_data2_reg_reg_15  ( .D(n6173), .CK(CLK), .Q(DOUT_47));
  QDFFHHD _i_CLEFIA128_data2_reg_reg_22  ( .D(n6180), .CK(CLK), .Q(DOUT_54));
  QDFFHHD _i_CLEFIA128_data2_reg_reg_14  ( .D(n6172), .CK(CLK), .Q(DOUT_46));
  QDFFHHD _i_CLEFIA128_data2_reg_reg_21  ( .D(n6179), .CK(CLK), .Q(DOUT_53));
  QDFFHHD _i_CLEFIA128_data2_reg_reg_13  ( .D(n6171), .CK(CLK), .Q(DOUT_45));
  QDFFHHD _i_CLEFIA128_data2_reg_reg_6  ( .D(n6164), .CK(CLK), .Q(DOUT_38));
  QDFFHHD _i_CLEFIA128_data2_reg_reg_4  ( .D(n6162), .CK(CLK), .Q(DOUT_36));
  QDFFHHD _i_CLEFIA128_data2_reg_reg_19  ( .D(n6177), .CK(CLK), .Q(DOUT_51));
  QDFFHHD _i_CLEFIA128_data2_reg_reg_17  ( .D(n6175), .CK(CLK), .Q(DOUT_49));
  QDFFHHD _i_CLEFIA128_data0_reg_reg_12  ( .D(n6202), .CK(CLK), .Q(DOUT_108));
  QDFFHHD _i_CLEFIA128_data0_reg_reg_29  ( .D(n6219), .CK(CLK), .Q(DOUT_125));
  QDFFHHD _i_CLEFIA128_data0_reg_reg_19  ( .D(n6209), .CK(CLK), .Q(DOUT_115));
  QDFFHHD _i_CLEFIA128_data2_reg_reg_10  ( .D(n6168), .CK(CLK), .Q(DOUT_42));
  QDFFHHD _i_CLEFIA128_data2_reg_reg_18  ( .D(n6176), .CK(CLK), .Q(DOUT_50));
  QDFFHHD _i_CLEFIA128_data2_reg_reg_11  ( .D(n6169), .CK(CLK), .Q(DOUT_43));
  QDFFHHD _i_CLEFIA128_data2_reg_reg_5  ( .D(n6163), .CK(CLK), .Q(DOUT_37));
  QDFFHHD _i_CLEFIA128_data2_reg_reg_1  ( .D(n6159), .CK(CLK), .Q(DOUT_33));
  QDFFHHD _i_CLEFIA128_data2_reg_reg_20  ( .D(n6178), .CK(CLK), .Q(DOUT_52));
  QDFFHHD _i_CLEFIA128_data2_reg_reg_3  ( .D(n6161), .CK(CLK), .Q(DOUT_35));
  QDFFHHD _i_CLEFIA128_data2_reg_reg_0  ( .D(n6221), .CK(CLK), .Q(DOUT_32));
  QDFFHHD _i_CLEFIA128_data3_reg_reg_0  ( .D(n6158), .CK(CLK), .Q(DOUT_0) );
  QDFFHHD _i_CLEFIA128_data2_reg_reg_25  ( .D(n6183), .CK(CLK), .Q(DOUT_57));
  QDFFHHD _i_CLEFIA128_data0_reg_reg_10  ( .D(n6200), .CK(CLK), .Q(DOUT_106));
  QDFFHHD _i_CLEFIA128_data0_reg_reg_20  ( .D(n6210), .CK(CLK), .Q(DOUT_116));
  QDFFHHD _i_CLEFIA128_data0_reg_reg_17  ( .D(n6207), .CK(CLK), .Q(DOUT_113));
  QDFFHHD _i_CLEFIA128_data0_reg_reg_25  ( .D(n6215), .CK(CLK), .Q(DOUT_121));
  QDFFHHD _i_CLEFIA128_data0_reg_reg_4  ( .D(n6194), .CK(CLK), .Q(DOUT_100));
  QDFFHHD _i_CLEFIA128_data1_reg_reg_4  ( .D(n6154), .CK(CLK), .Q(DOUT_68));
  QDFFHHD _i_CLEFIA128_data0_reg_reg_27  ( .D(n6217), .CK(CLK), .Q(DOUT_123));
  QDFFHHD _i_CLEFIA128_data0_reg_reg_30  ( .D(n6220), .CK(CLK), .Q(DOUT_126));
  QDFFHHD _i_CLEFIA128_data0_reg_reg_6  ( .D(n6196), .CK(CLK), .Q(DOUT_102));
  QDFFHHD _i_CLEFIA128_data0_reg_reg_31  ( .D(n6349), .CK(CLK), .Q(DOUT_127));
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_95  ( .D(n6254), .CK(CLK), .Q(_i_CLEFIA128_keyL _95) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_102  ( .D(n6247), .CK(CLK), .Q(_i_CLEFIA128_keyL _102) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_109  ( .D(n6240), .CK(CLK), .Q(_i_CLEFIA128_keyL _109) );
  QDFFHHD _i_CLEFIA128_data0_reg_reg_28  ( .D(n6218), .CK(CLK), .Q(DOUT_124));
  QDFFHHD _i_CLEFIA128_data0_reg_reg_21  ( .D(n6211), .CK(CLK), .Q(DOUT_117));
  QDFFHHD _i_CLEFIA128_data0_reg_reg_15  ( .D(n6205), .CK(CLK), .Q(DOUT_111));
  QDFFHHD _i_CLEFIA128_data0_reg_reg_23  ( .D(n6213), .CK(CLK), .Q(DOUT_119));
  QDFFHHD _i_CLEFIA128_data0_reg_reg_14  ( .D(n6204), .CK(CLK), .Q(DOUT_110));
  QDFFHHD _i_CLEFIA128_data0_reg_reg_5  ( .D(n6195), .CK(CLK), .Q(DOUT_101));
  QDFFHHD _i_CLEFIA128_data2_reg_reg_2  ( .D(n6160), .CK(CLK), .Q(DOUT_34));
  QDFFHHD _i_CLEFIA128_data3_reg_reg_2  ( .D(n6125), .CK(CLK), .Q(DOUT_2) );
  QDFFHHD _i_CLEFIA128_data0_reg_reg_2  ( .D(n6192), .CK(CLK), .Q(DOUT_98));
  QDFFHHD _i_CLEFIA128_data2_reg_reg_16  ( .D(n6174), .CK(CLK), .Q(DOUT_48));
  QDFFHHD _i_CLEFIA128_data1_reg_reg_16  ( .D(n6142), .CK(CLK), .Q(DOUT_80));
  QDFFHHD _i_CLEFIA128_data0_reg_reg_16  ( .D(n6206), .CK(CLK), .Q(DOUT_112));
  QDFFHHD _i_CLEFIA128_data2_reg_reg_9  ( .D(n6167), .CK(CLK), .Q(DOUT_41));
  QDFFHHD _i_CLEFIA128_data2_reg_reg_8  ( .D(n6166), .CK(CLK), .Q(DOUT_40));
  QDFFHHD _i_CLEFIA128_data1_reg_reg_8  ( .D(n6150), .CK(CLK), .Q(DOUT_72));
  QDFFHHD _i_CLEFIA128_data0_reg_reg_8  ( .D(n6198), .CK(CLK), .Q(DOUT_104));
  QDFFHHD _i_CLEFIA128_data0_reg_reg_3  ( .D(n6193), .CK(CLK), .Q(DOUT_99));
  QDFFHHD _i_CLEFIA128_data2_reg_reg_7  ( .D(n6165), .CK(CLK), .Q(DOUT_39));
  QDFFHHD _i_CLEFIA128_data3_reg_reg_7  ( .D(n6120), .CK(CLK), .Q(DOUT_7) );
  QDFFHHD _i_CLEFIA128_data0_reg_reg_7  ( .D(n6197), .CK(CLK), .Q(DOUT_103));
  QDFFHHD _i_CLEFIA128_data1_reg_reg_7  ( .D(n6151), .CK(CLK), .Q(DOUT_71));
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_88  ( .D(n6261), .CK(CLK), .Q(_i_CLEFIA128_keyL _88) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_81  ( .D(n6268), .CK(CLK), .Q(_i_CLEFIA128_keyL _81) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_74  ( .D(n6275), .CK(CLK), .Q(_i_CLEFIA128_keyL _74) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_67  ( .D(n6282), .CK(CLK), .Q(_i_CLEFIA128_keyL _67) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_123  ( .D(n6226), .CK(CLK), .Q(_i_CLEFIA128_keyL _123) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_116  ( .D(n6233), .CK(CLK), .Q(_i_CLEFIA128_keyL _116) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_17  ( .D(n6331), .CK(CLK), .Q(_i_CLEFIA128_keyL _17) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_24  ( .D(n6324), .CK(CLK), .Q(_i_CLEFIA128_keyL _24) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_31  ( .D(n6318), .CK(CLK), .Q(_i_CLEFIA128_keyL _31) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_38  ( .D(n6311), .CK(CLK), .Q(_i_CLEFIA128_keyL _38) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_45  ( .D(n6304), .CK(CLK), .Q(_i_CLEFIA128_keyL _45) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_52  ( .D(n6297), .CK(CLK), .Q(_i_CLEFIA128_keyL _52) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_59  ( .D(n6290), .CK(CLK), .Q(_i_CLEFIA128_keyL _59) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_3  ( .D(n6345), .CK(CLK), .Q(_i_CLEFIA128_keyL _3) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_10  ( .D(n6338), .CK(CLK), .Q(_i_CLEFIA128_keyL _10) );
  QDFFHHD _i_CLEFIA128_data0_reg_reg_24  ( .D(n6214), .CK(CLK), .Q(DOUT_120));
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_120  ( .D(n6229), .CK(CLK), .Q(_i_CLEFIA128_keyL _120) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_127  ( .D(n6222), .CK(CLK), .Q(_i_CLEFIA128_keyL _127) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_71  ( .D(n6278), .CK(CLK), .Q(_i_CLEFIA128_keyL _71) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_78  ( .D(n6271), .CK(CLK), .Q(_i_CLEFIA128_keyL _78) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_85  ( .D(n6264), .CK(CLK), .Q(_i_CLEFIA128_keyL _85) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_92  ( .D(n6257), .CK(CLK), .Q(_i_CLEFIA128_keyL _92) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_99  ( .D(n6250), .CK(CLK), .Q(_i_CLEFIA128_keyL _99) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_106  ( .D(n6243), .CK(CLK), .Q(_i_CLEFIA128_keyL _106) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_113  ( .D(n6236), .CK(CLK), .Q(_i_CLEFIA128_keyL _113) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_0  ( .D(n6348), .CK(CLK), .Q(_i_CLEFIA128_keyL _0) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_64  ( .D(n6285), .CK(CLK), .Q(_i_CLEFIA128_keyL _64) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_49  ( .D(n6300), .CK(CLK), .Q(_i_CLEFIA128_keyL _49) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_56  ( .D(n6293), .CK(CLK), .Q(_i_CLEFIA128_keyL _56) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_63  ( .D(n6286), .CK(CLK), .Q(_i_CLEFIA128_keyL _63) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_7  ( .D(n6341), .CK(CLK), .Q(_i_CLEFIA128_keyL _7) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_14  ( .D(n6334), .CK(CLK), .Q(_i_CLEFIA128_keyL _14) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_21  ( .D(n6327), .CK(CLK), .Q(_i_CLEFIA128_keyL _21) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_28  ( .D(n6350), .CK(CLK), .Q(_i_CLEFIA128_keyL _28) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_35  ( .D(n6314), .CK(CLK), .Q(_i_CLEFIA128_keyL _35) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_42  ( .D(n6307), .CK(CLK), .Q(_i_CLEFIA128_keyL _42) );
  QDFFHHD _i_CLEFIA128_data0_reg_reg_11  ( .D(n6201), .CK(CLK), .Q(DOUT_107));
  QDFFHHD _i_CLEFIA128_data1_reg_reg_11  ( .D(n6147), .CK(CLK), .Q(DOUT_75));
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_82  ( .D(n6267), .CK(CLK), .Q(_i_CLEFIA128_keyL _82) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_89  ( .D(n6260), .CK(CLK), .Q(_i_CLEFIA128_keyL _89) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_96  ( .D(n6253), .CK(CLK), .Q(_i_CLEFIA128_keyL _96) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_103  ( .D(n6246), .CK(CLK), .Q(_i_CLEFIA128_keyL _103) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_110  ( .D(n6239), .CK(CLK), .Q(_i_CLEFIA128_keyL _110) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_117  ( .D(n6232), .CK(CLK), .Q(_i_CLEFIA128_keyL _117) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_124  ( .D(n6225), .CK(CLK), .Q(_i_CLEFIA128_keyL _124) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_68  ( .D(n6281), .CK(CLK), .Q(_i_CLEFIA128_keyL _68) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_75  ( .D(n6274), .CK(CLK), .Q(_i_CLEFIA128_keyL _75) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_60  ( .D(n6289), .CK(CLK), .Q(_i_CLEFIA128_keyL _60) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_53  ( .D(n6296), .CK(CLK), .Q(_i_CLEFIA128_keyL _53) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_46  ( .D(n6303), .CK(CLK), .Q(_i_CLEFIA128_keyL _46) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_39  ( .D(n6310), .CK(CLK), .Q(_i_CLEFIA128_keyL _39) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_32  ( .D(n6317), .CK(CLK), .Q(_i_CLEFIA128_keyL _32) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_25  ( .D(n6323), .CK(CLK), .Q(_i_CLEFIA128_keyL _25) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_18  ( .D(n6330), .CK(CLK), .Q(_i_CLEFIA128_keyL _18) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_11  ( .D(n6337), .CK(CLK), .Q(_i_CLEFIA128_keyL _11) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_4  ( .D(n6344), .CK(CLK), .Q(_i_CLEFIA128_keyL _4) );
  QDFFHHD _i_CLEFIA128_data0_reg_reg_18  ( .D(n6208), .CK(CLK), .Q(DOUT_114));
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_77  ( .D(n6272), .CK(CLK), .Q(_i_CLEFIA128_keyL _77) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_84  ( .D(n6265), .CK(CLK), .Q(_i_CLEFIA128_keyL _84) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_91  ( .D(n6258), .CK(CLK), .Q(_i_CLEFIA128_keyL _91) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_98  ( .D(n6251), .CK(CLK), .Q(_i_CLEFIA128_keyL _98) );
  QDFFHHD _i_CLEFIA128_data0_reg_reg_1  ( .D(n6191), .CK(CLK), .Q(DOUT_97));
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_86  ( .D(n6263), .CK(CLK), .Q(_i_CLEFIA128_keyL _86) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_93  ( .D(n6256), .CK(CLK), .Q(_i_CLEFIA128_keyL _93) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_100  ( .D(n6249), .CK(CLK), .Q(_i_CLEFIA128_keyL _100) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_107  ( .D(n6242), .CK(CLK), .Q(_i_CLEFIA128_keyL _107) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_114  ( .D(n6235), .CK(CLK), .Q(_i_CLEFIA128_keyL _114) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_121  ( .D(n6228), .CK(CLK), .Q(_i_CLEFIA128_keyL _121) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_65  ( .D(n6284), .CK(CLK), .Q(_i_CLEFIA128_keyL _65) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_72  ( .D(n6277), .CK(CLK), .Q(_i_CLEFIA128_keyL _72) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_79  ( .D(n6270), .CK(CLK), .Q(_i_CLEFIA128_keyL _79) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_50  ( .D(n6299), .CK(CLK), .Q(_i_CLEFIA128_keyL _50) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_57  ( .D(n6292), .CK(CLK), .Q(_i_CLEFIA128_keyL _57) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_1  ( .D(n6347), .CK(CLK), .Q(_i_CLEFIA128_keyL _1) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_8  ( .D(n6340), .CK(CLK), .Q(_i_CLEFIA128_keyL _8) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_15  ( .D(n6333), .CK(CLK), .Q(_i_CLEFIA128_keyL _15) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_22  ( .D(n6326), .CK(CLK), .Q(_i_CLEFIA128_keyL _22) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_29  ( .D(n6320), .CK(CLK), .Q(_i_CLEFIA128_keyL _29) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_36  ( .D(n6313), .CK(CLK), .Q(_i_CLEFIA128_keyL _36) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_43  ( .D(n6306), .CK(CLK), .Q(_i_CLEFIA128_keyL _43) );
  QDFFHHD _i_CLEFIA128_data0_reg_reg_22  ( .D(n6212), .CK(CLK), .Q(DOUT_118));
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_118  ( .D(n6231), .CK(CLK), .Q(_i_CLEFIA128_keyL _118) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_125  ( .D(n6224), .CK(CLK), .Q(_i_CLEFIA128_keyL _125) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_69  ( .D(n6280), .CK(CLK), .Q(_i_CLEFIA128_keyL _69) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_76  ( .D(n6273), .CK(CLK), .Q(_i_CLEFIA128_keyL _76) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_83  ( .D(n6266), .CK(CLK), .Q(_i_CLEFIA128_keyL _83) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_90  ( .D(n6259), .CK(CLK), .Q(_i_CLEFIA128_keyL _90) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_97  ( .D(n6252), .CK(CLK), .Q(_i_CLEFIA128_keyL _97) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_104  ( .D(n6245), .CK(CLK), .Q(_i_CLEFIA128_keyL _104) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_111  ( .D(n6238), .CK(CLK), .Q(_i_CLEFIA128_keyL _111) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_26  ( .D(n6322), .CK(CLK), .Q(_i_CLEFIA128_keyL _26) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_33  ( .D(n6316), .CK(CLK), .Q(_i_CLEFIA128_keyL _33) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_40  ( .D(n6309), .CK(CLK), .Q(_i_CLEFIA128_keyL _40) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_47  ( .D(n6302), .CK(CLK), .Q(_i_CLEFIA128_keyL _47) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_54  ( .D(n6295), .CK(CLK), .Q(_i_CLEFIA128_keyL _54) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_61  ( .D(n6288), .CK(CLK), .Q(_i_CLEFIA128_keyL _61) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_5  ( .D(n6343), .CK(CLK), .Q(_i_CLEFIA128_keyL _5) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_12  ( .D(n6336), .CK(CLK), .Q(_i_CLEFIA128_keyL _12) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_19  ( .D(n6329), .CK(CLK), .Q(_i_CLEFIA128_keyL _19) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_73  ( .D(n6276), .CK(CLK), .Q(_i_CLEFIA128_keyL _73) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_80  ( .D(n6269), .CK(CLK), .Q(_i_CLEFIA128_keyL _80) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_87  ( .D(n6262), .CK(CLK), .Q(_i_CLEFIA128_keyL _87) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_94  ( .D(n6255), .CK(CLK), .Q(_i_CLEFIA128_keyL _94) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_101  ( .D(n6248), .CK(CLK), .Q(_i_CLEFIA128_keyL _101) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_108  ( .D(n6241), .CK(CLK), .Q(_i_CLEFIA128_keyL _108) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_115  ( .D(n6234), .CK(CLK), .Q(_i_CLEFIA128_keyL _115) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_122  ( .D(n6227), .CK(CLK), .Q(_i_CLEFIA128_keyL _122) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_66  ( .D(n6283), .CK(CLK), .Q(_i_CLEFIA128_keyL _66) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_51  ( .D(n6298), .CK(CLK), .Q(_i_CLEFIA128_keyL _51) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_58  ( .D(n6291), .CK(CLK), .Q(_i_CLEFIA128_keyL _58) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_2  ( .D(n6346), .CK(CLK), .Q(_i_CLEFIA128_keyL _2) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_9  ( .D(n6339), .CK(CLK), .Q(_i_CLEFIA128_keyL _9) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_16  ( .D(n6332), .CK(CLK), .Q(_i_CLEFIA128_keyL _16) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_23  ( .D(n6325), .CK(CLK), .Q(_i_CLEFIA128_keyL _23) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_30  ( .D(n6319), .CK(CLK), .Q(_i_CLEFIA128_keyL _30) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_37  ( .D(n6312), .CK(CLK), .Q(_i_CLEFIA128_keyL _37) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_44  ( .D(n6305), .CK(CLK), .Q(_i_CLEFIA128_keyL _44) );
  QDFFHHD _i_CLEFIA128_data0_reg_reg_9  ( .D(n6199), .CK(CLK), .Q(DOUT_105));
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_105  ( .D(n6244), .CK(CLK), .Q(_i_CLEFIA128_keyL _105) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_112  ( .D(n6237), .CK(CLK), .Q(_i_CLEFIA128_keyL _112) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_119  ( .D(n6230), .CK(CLK), .Q(_i_CLEFIA128_keyL _119) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_126  ( .D(n6223), .CK(CLK), .Q(_i_CLEFIA128_keyL _126) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_70  ( .D(n6279), .CK(CLK), .Q(_i_CLEFIA128_keyL _70) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_55  ( .D(n6294), .CK(CLK), .Q(_i_CLEFIA128_keyL _55) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_62  ( .D(n6287), .CK(CLK), .Q(_i_CLEFIA128_keyL _62) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_6  ( .D(n6342), .CK(CLK), .Q(_i_CLEFIA128_keyL _6) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_13  ( .D(n6335), .CK(CLK), .Q(_i_CLEFIA128_keyL _13) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_20  ( .D(n6328), .CK(CLK), .Q(_i_CLEFIA128_keyL _20) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_27  ( .D(n6321), .CK(CLK), .Q(_i_CLEFIA128_keyL _27) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_34  ( .D(n6315), .CK(CLK), .Q(_i_CLEFIA128_keyL _34) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_41  ( .D(n6308), .CK(CLK), .Q(_i_CLEFIA128_keyL _41) );
  QDFFHHD _i_CLEFIA128_keyL_reg_reg_48  ( .D(n6301), .CK(CLK), .Q(_i_CLEFIA128_keyL _48) );
  QDFFHHD _i_CLEFIA128_data1_reg_reg_9  ( .D(n6149), .CK(CLK), .Q(DOUT_73));
  QDFFHHD _i_CLEFIA128_data1_reg_reg_22  ( .D(n6136), .CK(CLK), .Q(DOUT_86));
  QDFFHHD _i_CLEFIA128_data1_reg_reg_1  ( .D(n6157), .CK(CLK), .Q(DOUT_65));
  QDFFHHD _i_CLEFIA128_data0_reg_reg_13  ( .D(n6203), .CK(CLK), .Q(DOUT_109));
  QDFFHHD _i_CLEFIA128_data1_reg_reg_13  ( .D(n6145), .CK(CLK), .Q(DOUT_77));
  QDFFHHD _i_CLEFIA128_data1_reg_reg_18  ( .D(n6140), .CK(CLK), .Q(DOUT_82));
  QDFFHHD _i_CLEFIA128_data1_reg_reg_24  ( .D(n6134), .CK(CLK), .Q(DOUT_88));
  QDFFHHD _i_CLEFIA128_data1_reg_reg_3  ( .D(n6155), .CK(CLK), .Q(DOUT_67));
  QDFFHHD _i_CLEFIA128_data3_reg_reg_8  ( .D(n6119), .CK(CLK), .Q(DOUT_8) );
  QDFFHHD _i_CLEFIA128_data3_reg_reg_9  ( .D(n6118), .CK(CLK), .Q(DOUT_9) );
  QDFFHHD _i_CLEFIA128_data3_reg_reg_16  ( .D(n6111), .CK(CLK), .Q(DOUT_16));
  QDFFHHD _i_CLEFIA128_data1_reg_reg_2  ( .D(n6156), .CK(CLK), .Q(DOUT_66));
  QDFFHHD _i_CLEFIA128_data1_reg_reg_5  ( .D(n6153), .CK(CLK), .Q(DOUT_69));
  QDFFHHD _i_CLEFIA128_data1_reg_reg_14  ( .D(n6144), .CK(CLK), .Q(DOUT_78));
  QDFFHHD _i_CLEFIA128_data1_reg_reg_23  ( .D(n6135), .CK(CLK), .Q(DOUT_87));
  QDFFHHD _i_CLEFIA128_data1_reg_reg_15  ( .D(n6143), .CK(CLK), .Q(DOUT_79));
  QDFFHHD _i_CLEFIA128_data1_reg_reg_21  ( .D(n6137), .CK(CLK), .Q(DOUT_85));
  QDFFHHD _i_CLEFIA128_data1_reg_reg_28  ( .D(n6130), .CK(CLK), .Q(DOUT_92));
  QDFFHHD _i_CLEFIA128_data1_reg_reg_31  ( .D(n6127), .CK(CLK), .Q(DOUT_95));
  QDFFHHD _i_CLEFIA128_data1_reg_reg_6  ( .D(n6152), .CK(CLK), .Q(DOUT_70));
  QDFFHHD _i_CLEFIA128_data1_reg_reg_30  ( .D(n6128), .CK(CLK), .Q(DOUT_94));
  QDFFHHD _i_CLEFIA128_data1_reg_reg_27  ( .D(n6131), .CK(CLK), .Q(DOUT_91));
  QDFFHHD _i_CLEFIA128_data1_reg_reg_25  ( .D(n6133), .CK(CLK), .Q(DOUT_89));
  QDFFHHD _i_CLEFIA128_data1_reg_reg_17  ( .D(n6141), .CK(CLK), .Q(DOUT_81));
  QDFFHHD _i_CLEFIA128_data1_reg_reg_20  ( .D(n6138), .CK(CLK), .Q(DOUT_84));
  QDFFHHD _i_CLEFIA128_data3_reg_reg_10  ( .D(n6117), .CK(CLK), .Q(DOUT_10));
  QDFFHHD _i_CLEFIA128_data3_reg_reg_25  ( .D(n6102), .CK(CLK), .Q(DOUT_25));
  QDFFHHD _i_CLEFIA128_data3_reg_reg_3  ( .D(n6124), .CK(CLK), .Q(DOUT_3) );
  QDFFHHD _i_CLEFIA128_data3_reg_reg_20  ( .D(n6107), .CK(CLK), .Q(DOUT_20));
  QDFFHHD _i_CLEFIA128_data3_reg_reg_1  ( .D(n6126), .CK(CLK), .Q(DOUT_1) );
  QDFFHHD _i_CLEFIA128_data3_reg_reg_5  ( .D(n6122), .CK(CLK), .Q(DOUT_5) );
  QDFFHHD _i_CLEFIA128_data3_reg_reg_11  ( .D(n6116), .CK(CLK), .Q(DOUT_11));
  QDFFHHD _i_CLEFIA128_data3_reg_reg_18  ( .D(n6109), .CK(CLK), .Q(DOUT_18));
  QDFFHHD _i_CLEFIA128_data1_reg_reg_10  ( .D(n6148), .CK(CLK), .Q(DOUT_74));
  QDFFHHD _i_CLEFIA128_data1_reg_reg_19  ( .D(n6139), .CK(CLK), .Q(DOUT_83));
  QDFFHHD _i_CLEFIA128_data1_reg_reg_29  ( .D(n6129), .CK(CLK), .Q(DOUT_93));
  QDFFHHD _i_CLEFIA128_data3_reg_reg_12  ( .D(n6115), .CK(CLK), .Q(DOUT_12));
  QDFFHHD _i_CLEFIA128_data3_reg_reg_17  ( .D(n6110), .CK(CLK), .Q(DOUT_17));
  QDFFHHD _i_CLEFIA128_data3_reg_reg_19  ( .D(n6108), .CK(CLK), .Q(DOUT_19));
  QDFFHHD _i_CLEFIA128_data3_reg_reg_4  ( .D(n6123), .CK(CLK), .Q(DOUT_4) );
  QDFFHHD _i_CLEFIA128_data3_reg_reg_6  ( .D(n6121), .CK(CLK), .Q(DOUT_6) );
  QDFFHHD _i_CLEFIA128_data3_reg_reg_13  ( .D(n6114), .CK(CLK), .Q(DOUT_13));
  QDFFHHD _i_CLEFIA128_data3_reg_reg_21  ( .D(n6106), .CK(CLK), .Q(DOUT_21));
  QDFFHHD _i_CLEFIA128_data3_reg_reg_14  ( .D(n6113), .CK(CLK), .Q(DOUT_14));
  QDFFHHD _i_CLEFIA128_data3_reg_reg_22  ( .D(n6105), .CK(CLK), .Q(DOUT_22));
  QDFFHHD _i_CLEFIA128_data3_reg_reg_15  ( .D(n6112), .CK(CLK), .Q(DOUT_15));
  QDFFHHD _i_CLEFIA128_data3_reg_reg_23  ( .D(n6104), .CK(CLK), .Q(DOUT_23));
  QDFFHHD _i_CLEFIA128_data1_reg_reg_12  ( .D(n6146), .CK(CLK), .Q(DOUT_76));
  QDFFHHD _i_CLEFIA128_data3_reg_reg_26  ( .D(n6101), .CK(CLK), .Q(DOUT_26));
  QDFFHHD _i_CLEFIA128_data3_reg_reg_28  ( .D(n6099), .CK(CLK), .Q(DOUT_28));
  QDFFHHD _i_CLEFIA128_data3_reg_reg_27  ( .D(n6100), .CK(CLK), .Q(DOUT_27));
  QDFFHHD _i_CLEFIA128_data3_reg_reg_24  ( .D(n6103), .CK(CLK), .Q(DOUT_24));
  QDFFHHD _i_CLEFIA128_data3_reg_reg_29  ( .D(n6098), .CK(CLK), .Q(DOUT_29));
  QDFFHHD _i_CLEFIA128_data3_reg_reg_30  ( .D(n6097), .CK(CLK), .Q(DOUT_30));
  QDFFHHD _i_CLEFIA128_data3_reg_reg_31  ( .D(n6096), .CK(CLK), .Q(DOUT_31));
  QDFFHHD _i_CLEFIA128_data1_reg_reg_26  ( .D(n6132), .CK(CLK), .Q(DOUT_90));
  DFFHHD _i_CLEFIA128_rndcnt_reg_reg_1  ( .D(n6370), .CK(CLK), .Q(n8797), .QB(n8798) );
  DFCRBEHD _i_CLEFIA128_DVLD_reg_reg  ( .D(n15523), .RB(n15522), .CK(CLK), .Q(DVLD), .QB(n15521) );
  ND2CHD U6504 ( .I1(n15095), .I2(n7043), .O(n7352) );
  ND2HHD U6505 ( .I1(n9867), .I2(n15500), .O(n10192) );
  ND2DHD U6506 ( .I1(n15235), .I2(n15500), .O(n8090) );
  ND2DHD U6507 ( .I1(n15024), .I2(n11130), .O(n7210) );
  ND2DHD U6508 ( .I1(n15207), .I2(n14786), .O(n14794) );
  MUX2EHD U6509 ( .A(n13733), .B(n13732), .S(n14573), .O(n9141) );
  ND2DHD U6510 ( .I1(n15440), .I2(n8277), .O(n9767) );
  MUX2EHD U6511 ( .A(n13781), .B(n13780), .S(n15374), .O(n13789) );
  ND2DHD U6512 ( .I1(n15171), .I2(n15500), .O(n7901) );
  ND2DHD U6513 ( .I1(n8011), .I2(n15311), .O(n8010) );
  ND2HHD U6514 ( .I1(n9867), .I2(n11130), .O(n9328) );
  ND2HHD U6515 ( .I1(n7952), .I2(n11130), .O(n6638) );
  AOI22BHD U6516 ( .A1(n7045), .A2(n14285), .B1(n15504), .B2(n14284), .O(n14286) );
  ND2DHD U6517 ( .I1(n14647), .I2(n13927), .O(n7111) );
  ND2DHD U6518 ( .I1(n15095), .I2(n15500), .O(n14110) );
  AN2EHD U6519 ( .I1(n8602), .I2(n13965), .O(n8601) );
  BUFJHD U6520 ( .I(n15439), .O(n6604) );
  ND2DHD U6521 ( .I1(n14938), .I2(n8287), .O(n10197) );
  OR2HHD U6522 ( .I1(n15450), .I2(n15449), .O(n15454) );
  NR2GHD U6523 ( .I1(n8313), .I2(n9109), .O(n9108) );
  NR2GHD U6524 ( .I1(n14348), .I2(n14347), .O(n7135) );
  NR2CHD U6525 ( .I1(n13047), .I2(n13046), .O(n13048) );
  NR2CHD U6526 ( .I1(n12823), .I2(n12822), .O(n12824) );
  NR2CHD U6527 ( .I1(n14254), .I2(n14253), .O(n14255) );
  AO22CHD U6528 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _115), .B1(n15504), .B2(_i_CLEFIA128_keyK _51), .O(n8284) );
  INVDHD U6529 ( .I(n15513), .O(n6556) );
  INVGHD U6530 ( .I(n15307), .O(n8705) );
  AO22CHD U6531 ( .A1(n8121), .A2(n7045), .B1(n15504), .B2(n13041), .O(n8451));
  XNR2HHD U6532 ( .I1(n8068), .I2(n8067), .O(n8011) );
  INVJHD U6533 ( .I(n8468), .O(n8466) );
  AO22CHD U6534 ( .A1(n7045), .A2(n14296), .B1(n15504), .B2(n14295), .O(n8258));
  AO22CHD U6535 ( .A1(n7045), .A2(n14350), .B1(n15504), .B2(n14349), .O(n8261));
  AO22CHD U6536 ( .A1(n7045), .A2(n15217), .B1(n15504), .B2(n15216), .O(n15218) );
  ND2HHD U6537 ( .I1(n14465), .I2(_i_CLEFIA128_CON_T_x _1), .O(n14738) );
  NR2GHD U6538 ( .I1(n12887), .I2(n7186), .O(n8877) );
  BUFHHD U6539 ( .I(n14705), .O(n9538) );
  XNR2CHD U6540 ( .I1(DIN_67), .I2(_i_CLEFIA128_keyK _99), .O(n14337) );
  XOR2EHD U6541 ( .I1(n8761), .I2(n8870), .O(n7214) );
  XNR2EHD U6542 ( .I1(n14108), .I2(n9776), .O(n7175) );
  XOR2EHD U6543 ( .I1(DOUT_16), .I2(n9797), .O(n13779) );
  INVGHD U6544 ( .I(_i_CLEFIA128_keyL _117), .O(n14943) );
  INVGHD U6545 ( .I(_i_CLEFIA128_keyL _61), .O(n15285) );
  INVCHD U6546 ( .I(_i_CLEFIA128_keyK _99), .O(n14326) );
  BUFDHD U6547 ( .I(n6724), .O(n7048) );
  INVDHD U6548 ( .I(_i_CLEFIA128_CON_T_x _1), .O(n14464) );
  XOR2EHD U6549 ( .I1(n7607), .I2(n6847), .O(n14014) );
  INVDHD U6550 ( .I(n9768), .O(n9409) );
  XOR2EHD U6551 ( .I1(n7195), .I2(n14169), .O(n14493) );
  XOR2EHD U6552 ( .I1(n14028), .I2(n6852), .O(n14005) );
  INVDHD U6553 ( .I(_i_CLEFIA128_keyL _22), .O(n15201) );
  INVDHD U6554 ( .I(_i_CLEFIA128_keyL _109), .O(n14483) );
  XNR2EHD U6555 ( .I1(n8561), .I2(n13715), .O(n13895) );
  BUFIHD U6556 ( .I(n14329), .O(n9775) );
  XOR2EHD U6557 ( .I1(n9761), .I2(n8756), .O(n13912) );
  XNR2EHD U6558 ( .I1(n14330), .I2(n14634), .O(n14333) );
  BUFHHD U6559 ( .I(n8309), .O(n6889) );
  BUFCKHHD U6560 ( .I(n13717), .O(n9657) );
  XOR2EHD U6561 ( .I1(n7832), .I2(n14106), .O(n7506) );
  XNR2EHD U6562 ( .I1(n14168), .I2(n6808), .O(n8418) );
  XNR2EHD U6563 ( .I1(DOUT_74), .I2(n7836), .O(n7572) );
  XNR2CHD U6564 ( .I1(DOUT_78), .I2(n14028), .O(n14029) );
  INVDHD U6565 ( .I(n10160), .O(n8761) );
  XOR2EHD U6566 ( .I1(n8064), .I2(n14215), .O(n8063) );
  BUFJHD U6567 ( .I(n14994), .O(n8870) );
  XOR2EHD U6568 ( .I1(DOUT_30), .I2(n9757), .O(n9024) );
  BUFHHD U6569 ( .I(n7607), .O(n7110) );
  INVGHD U6570 ( .I(n14636), .O(n10019) );
  BUFIHD U6571 ( .I(n6874), .O(n9768) );
  XNR2HHD U6572 ( .I1(n9664), .I2(n14028), .O(n14213) );
  BUFHHD U6573 ( .I(n10149), .O(n7932) );
  BUFKHD U6574 ( .I(n13951), .O(n9960) );
  ND2HHD U6575 ( .I1(n13850), .I2(n13851), .O(n14215) );
  INVCHD U6576 ( .I(ENCDEC), .O(n10911) );
  ND2HHD U6577 ( .I1(n7080), .I2(n13052), .O(n14227) );
  ND2HHD U6578 ( .I1(n10923), .I2(n10922), .O(n15450) );
  ND2DHD U6579 ( .I1(n14407), .I2(n14403), .O(n14709) );
  OR2EHD U6580 ( .I1(n14678), .I2(n14683), .O(n10300) );
  INVCHD U6581 ( .I(DOUT_94), .O(n7832) );
  BUFJHD U6582 ( .I(n14138), .O(n9013) );
  ND2CHD U6583 ( .I1(n14688), .I2(_i_CLEFIA128_state_reg _1), .O(n10923) );
  INVJHD U6584 ( .I(n6739), .O(n6808) );
  AN2CHD U6585 ( .I1(n14444), .I2(BSY), .O(n10922) );
  BUFIHD U6586 ( .I(n8790), .O(n6577) );
  XNR2CHD U6587 ( .I1(DOUT_11), .I2(n7100), .O(n6800) );
  NR2EHD U6588 ( .I1(n13555), .I2(n13554), .O(n7945) );
  NR2CHD U6589 ( .I1(n14678), .I2(n14685), .O(n10302) );
  INVDHD U6590 ( .I(SRST), .O(n14430) );
  OA13EHD U6591 ( .B1(n13658), .B2(n13657), .B3(n13848), .A1(n13835), .O(n13669) );
  INVHHD U6592 ( .I(n6636), .O(n8788) );
  INVHHD U6593 ( .I(n14167), .O(n9415) );
  INVDHD U6594 ( .I(DOUT_92), .O(n9496) );
  INVJHD U6595 ( .I(n7813), .O(n8309) );
  INVJHD U6596 ( .I(n7357), .O(n8030) );
  NR2EHD U6597 ( .I1(n12085), .I2(n12084), .O(n9805) );
  INVGHD U6598 ( .I(n13111), .O(n13109) );
  NR2EHD U6599 ( .I1(n9537), .I2(n13112), .O(n9536) );
  INVLHD U6600 ( .I(n7916), .O(n7917) );
  AN2CHD U6601 ( .I1(n9378), .I2(n12842), .O(n9377) );
  INVCHD U6602 ( .I(n10105), .O(n7405) );
  AN2EHD U6603 ( .I1(n11211), .I2(n11230), .O(n9683) );
  ND3CHD U6604 ( .I1(n7508), .I2(n11231), .I3(n10635), .O(n10683) );
  ND2DHD U6605 ( .I1(n12548), .I2(n12646), .O(n12549) );
  ND3CHD U6606 ( .I1(n7179), .I2(n10288), .I3(n10287), .O(n10286) );
  ND3CHD U6607 ( .I1(n13650), .I2(n13649), .I3(n8242), .O(n13658) );
  ND2CHD U6608 ( .I1(n13621), .I2(n13193), .O(n13206) );
  ND2HHD U6609 ( .I1(n7602), .I2(n11216), .O(n7601) );
  NR2BHD U6610 ( .I1(n10129), .I2(n12122), .O(n13168) );
  INVDHD U6611 ( .I(n6855), .O(n6790) );
  INVGHD U6612 ( .I(BSY), .O(n14678) );
  INVCHD U6613 ( .I(n10792), .O(n10667) );
  INVDHD U6614 ( .I(n12492), .O(n10277) );
  INVCHD U6615 ( .I(n12752), .O(n6611) );
  NR2BHD U6616 ( .I1(n13679), .I2(n8582), .O(n13509) );
  NR2EHD U6617 ( .I1(n14069), .I2(n13245), .O(n13250) );
  BUFIHD U6618 ( .I(n8624), .O(n6533) );
  ND3CHD U6619 ( .I1(n13213), .I2(n13211), .I3(n13212), .O(n13214) );
  NR2EHD U6620 ( .I1(n13495), .I2(n7764), .O(n9508) );
  NR2EHD U6621 ( .I1(n11215), .I2(n9331), .O(n7834) );
  AN2CHD U6622 ( .I1(n13179), .I2(n13178), .O(n8712) );
  BUFCKHHD U6623 ( .I(n13636), .O(n9878) );
  INVCHD U6624 ( .I(n13141), .O(n6507) );
  NR2EHD U6625 ( .I1(n13032), .I2(n8672), .O(n8671) );
  AN2EHD U6626 ( .I1(n8654), .I2(n13819), .O(n8395) );
  NR3BHD U6627 ( .I1(n11414), .I2(n10514), .I3(n11409), .O(n6793) );
  NR2EHD U6628 ( .I1(n10125), .I2(n13368), .O(n13369) );
  NR2EHD U6629 ( .I1(n13202), .I2(n13201), .O(n13203) );
  NR2CHD U6630 ( .I1(n12249), .I2(n12250), .O(n8670) );
  INVDHD U6631 ( .I(n13181), .O(n8711) );
  ND3CHD U6632 ( .I1(n9740), .I2(n7019), .I3(n10035), .O(n9071) );
  ND3CHD U6633 ( .I1(n13391), .I2(n13390), .I3(n13389), .O(n13392) );
  ND2DHD U6634 ( .I1(n9241), .I2(n9240), .O(n12072) );
  ND2HHD U6635 ( .I1(n6978), .I2(n8563), .O(n8949) );
  NR2BHD U6636 ( .I1(n8846), .I2(n13523), .O(n13529) );
  ND2CHD U6637 ( .I1(n8652), .I2(n9405), .O(n8619) );
  ND2DHD U6638 ( .I1(n13278), .I2(n10299), .O(n14683) );
  NR2CHD U6639 ( .I1(n14069), .I2(n14068), .O(n7714) );
  ND2DHD U6640 ( .I1(n9468), .I2(n9466), .O(n12838) );
  NR2EHD U6641 ( .I1(n8580), .I2(n12845), .O(n12855) );
  INVDHD U6642 ( .I(n13622), .O(n13141) );
  INVDHD U6643 ( .I(n9236), .O(n9240) );
  INVGHD U6644 ( .I(n12672), .O(n8580) );
  ND2DHD U6645 ( .I1(n9123), .I2(n9221), .O(n9122) );
  OA12EHD U6646 ( .B1(n12055), .B2(n13169), .A1(n13585), .O(n6555) );
  INVHHD U6647 ( .I(n13095), .O(n14066) );
  NR2CHD U6648 ( .I1(n9454), .I2(n9467), .O(n9466) );
  INVDHD U6649 ( .I(n12978), .O(n8672) );
  OR3EHD U6650 ( .I1(n12496), .I2(n11435), .I3(n9388), .O(n10993) );
  INVCHD U6651 ( .I(n7441), .O(n13390) );
  NR2EHD U6652 ( .I1(n9182), .I2(n14057), .O(n9181) );
  INVDHD U6653 ( .I(n12746), .O(n8682) );
  AN2EHD U6654 ( .I1(n12454), .I2(n12456), .O(n11187) );
  NR2EHD U6655 ( .I1(n13836), .I2(n12090), .O(n9405) );
  NR2EHD U6656 ( .I1(n12070), .I2(n12071), .O(n9241) );
  NR2EHD U6657 ( .I1(n11157), .I2(n11447), .O(n9088) );
  ND3CHD U6658 ( .I1(n10989), .I2(n6858), .I3(n10988), .O(n10994) );
  NR2EHD U6659 ( .I1(n11373), .I2(n11372), .O(n11374) );
  NR2EHD U6660 ( .I1(n7273), .I2(n7271), .O(n7270) );
  NR2EHD U6661 ( .I1(n8003), .I2(n8002), .O(n11344) );
  NR2EHD U6662 ( .I1(n7847), .I2(n7562), .O(n7561) );
  NR2BHD U6663 ( .I1(n8595), .I2(n14045), .O(n9403) );
  NR2CHD U6664 ( .I1(n11136), .I2(n11137), .O(n8906) );
  ND3CHD U6665 ( .I1(n13057), .I2(n13056), .I3(n13055), .O(n13065) );
  AN2EHD U6666 ( .I1(n12093), .I2(n9154), .O(n12094) );
  ND2DHD U6667 ( .I1(n13063), .I2(n13062), .O(n13498) );
  OR3EHD U6668 ( .I1(n13244), .I2(n13236), .I3(n13235), .O(n13237) );
  ND3CHD U6669 ( .I1(n11493), .I2(n11492), .I3(n12555), .O(n11502) );
  NR2CHD U6670 ( .I1(n12232), .I2(n12231), .O(n12236) );
  NR2CHD U6671 ( .I1(n10103), .I2(n10104), .O(n10102) );
  ND2CHD U6672 ( .I1(n11220), .I2(n8785), .O(n10047) );
  ND3CHD U6673 ( .I1(n12456), .I2(n12455), .I3(n8781), .O(n12460) );
  OR3EHD U6674 ( .I1(n12528), .I2(n12530), .I3(n12529), .O(n12531) );
  NR2CHD U6675 ( .I1(n8770), .I2(n7899), .O(n11151) );
  BUFIHD U6676 ( .I(n13170), .O(n9629) );
  ND3CHD U6677 ( .I1(n6514), .I2(n13038), .I3(n9245), .O(n9243) );
  ND2DHD U6678 ( .I1(n8416), .I2(n9646), .O(n8057) );
  ND3CHD U6679 ( .I1(n10433), .I2(n10432), .I3(n10434), .O(n8527) );
  OR3CHD U6680 ( .I1(n11725), .I2(n13647), .I3(n11724), .O(n11729) );
  INVDHD U6681 ( .I(_i_CLEFIA128_rndcnt_reg _3), .O(n14415) );
  NR2CHD U6682 ( .I1(n7264), .I2(n11050), .O(n11051) );
  NR2BHD U6683 ( .I1(n13584), .I2(n13117), .O(n13118) );
  AN3EHD U6684 ( .I1(n10696), .I2(n12464), .I3(n9034), .O(n7898) );
  NR2CHD U6685 ( .I1(n10765), .I2(n10892), .O(n8493) );
  AN2CHD U6686 ( .I1(n13208), .I2(n13183), .O(n13142) );
  AN3EHD U6687 ( .I1(n10850), .I2(n7606), .I3(n7375), .O(n10360) );
  AN2EHD U6688 ( .I1(n9709), .I2(n12518), .O(n12519) );
  INVHHD U6689 ( .I(n8828), .O(n6705) );
  INVDHD U6690 ( .I(n12503), .O(n10251) );
  INVCHD U6691 ( .I(n8919), .O(n10453) );
  AN2EHD U6692 ( .I1(n9224), .I2(n12451), .O(n11287) );
  INVDHD U6693 ( .I(n11212), .O(n11214) );
  AN2CHD U6694 ( .I1(n12454), .I2(n12464), .O(n8426) );
  INVDHD U6695 ( .I(n9492), .O(n9486) );
  NR2EHD U6696 ( .I1(n11448), .I2(n9196), .O(n9195) );
  ND3CHD U6697 ( .I1(n13844), .I2(n13512), .I3(n13804), .O(n9001) );
  BUFCKIHD U6698 ( .I(n9742), .O(n7077) );
  NR2EHD U6699 ( .I1(n10595), .I2(n11177), .O(n10597) );
  NR2EHD U6700 ( .I1(n13834), .I2(n7418), .O(n7926) );
  ND2DHD U6701 ( .I1(n12747), .I2(n12768), .O(n11044) );
  AN2CHD U6702 ( .I1(n6753), .I2(n9398), .O(n12248) );
  AN3EHD U6703 ( .I1(n11644), .I2(n13099), .I3(n10296), .O(n14047) );
  AN3EHD U6704 ( .I1(n7382), .I2(n6535), .I3(n10080), .O(n12924) );
  AN3EHD U6705 ( .I1(n12265), .I2(n9770), .I3(n13589), .O(n12923) );
  INVGHD U6706 ( .I(n7593), .O(n12200) );
  NR2EHD U6707 ( .I1(n11494), .I2(n11495), .O(n11499) );
  NR2EHD U6708 ( .I1(n11394), .I2(n11395), .O(n12776) );
  INVDHD U6709 ( .I(n7396), .O(n9713) );
  INVGHD U6710 ( .I(n12565), .O(n7660) );
  INVCHD U6711 ( .I(n13235), .O(n13069) );
  NR2EHD U6712 ( .I1(n10649), .I2(n10650), .O(n7364) );
  NR2EHD U6713 ( .I1(n13682), .I2(n8818), .O(n13531) );
  BUFCKHHD U6714 ( .I(n14080), .O(n6707) );
  INVDHD U6715 ( .I(n12211), .O(n13229) );
  NR2EHD U6716 ( .I1(n11101), .I2(n11102), .O(n11377) );
  INVDHD U6717 ( .I(n6515), .O(n6514) );
  INVDHD U6718 ( .I(n12716), .O(n9326) );
  AN2EHD U6719 ( .I1(n8832), .I2(n13506), .O(n13661) );
  ND2CHD U6720 ( .I1(n6682), .I2(n13844), .O(n13524) );
  NR2EHD U6721 ( .I1(n13082), .I2(n13081), .O(n14075) );
  NR2EHD U6722 ( .I1(n12345), .I2(n12344), .O(n13429) );
  NR2EHD U6723 ( .I1(n13235), .I2(n13054), .O(n13056) );
  NR2EHD U6724 ( .I1(n13129), .I2(n10013), .O(n13601) );
  NR2EHD U6725 ( .I1(n8491), .I2(n9382), .O(n8490) );
  ND2HHD U6726 ( .I1(n8350), .I2(n9146), .O(n6813) );
  NR2EHD U6727 ( .I1(n7445), .I2(n7446), .O(n7084) );
  BUFHHD U6728 ( .I(n13681), .O(n9094) );
  INVGHD U6729 ( .I(n6888), .O(n12545) );
  OR2EHD U6730 ( .I1(n9299), .I2(n11708), .O(n9068) );
  NR2EHD U6731 ( .I1(n11141), .I2(n9446), .O(n11146) );
  NR2EHD U6732 ( .I1(n11131), .I2(n11132), .O(n11133) );
  NR2EHD U6733 ( .I1(n10359), .I2(n10358), .O(n10361) );
  BUFGHD U6734 ( .I(n12211), .O(n8993) );
  INVJHD U6735 ( .I(n11651), .O(n11822) );
  NR2EHD U6736 ( .I1(n8673), .I2(n8322), .O(n12978) );
  NR2EHD U6737 ( .I1(n12680), .I2(n12679), .O(n7818) );
  NR2EHD U6738 ( .I1(n7493), .I2(n7492), .O(n7495) );
  NR2EHD U6739 ( .I1(n12860), .I2(n12813), .O(n9379) );
  NR2EHD U6740 ( .I1(n7448), .I2(n7447), .O(n7444) );
  BUFHHD U6741 ( .I(n10892), .O(n7793) );
  AN2HHD U6742 ( .I1(n11312), .I2(n10628), .O(n12474) );
  NR2EHD U6743 ( .I1(n7665), .I2(n11405), .O(n7659) );
  NR2EHD U6744 ( .I1(n11486), .I2(n9600), .O(n10064) );
  INVDHD U6745 ( .I(n11272), .O(n7913) );
  INVJHD U6746 ( .I(n12576), .O(n6568) );
  NR2GHD U6747 ( .I1(n10067), .I2(n9795), .O(n12590) );
  NR2EHD U6748 ( .I1(n9662), .I2(n11731), .O(n9542) );
  NR2EHD U6749 ( .I1(n10221), .I2(n6549), .O(n8432) );
  NR2EHD U6750 ( .I1(n9081), .I2(n13017), .O(n9121) );
  NR2EHD U6751 ( .I1(n12505), .I2(n12494), .O(n10987) );
  INVGHD U6752 ( .I(n8823), .O(n10707) );
  NR2EHD U6753 ( .I1(n11473), .I2(n11474), .O(n11478) );
  AN2EHD U6754 ( .I1(n7701), .I2(n13833), .O(n8857) );
  NR2EHD U6755 ( .I1(n12744), .I2(n8869), .O(n7710) );
  AN2HHD U6756 ( .I1(n12054), .I2(n12062), .O(n13622) );
  INVDHD U6757 ( .I(n12054), .O(n12063) );
  OR2CHD U6758 ( .I1(n9441), .I2(n10809), .O(n8421) );
  NR2EHD U6759 ( .I1(n8453), .I2(n11487), .O(n10065) );
  ND2DHD U6760 ( .I1(n8365), .I2(n10282), .O(n8952) );
  ND2HHD U6761 ( .I1(n11636), .I2(n14079), .O(n13075) );
  NR2CHD U6762 ( .I1(n9434), .I2(n13825), .O(n9432) );
  AN2EHD U6763 ( .I1(n11318), .I2(n11300), .O(n12506) );
  NR2EHD U6764 ( .I1(n11183), .I2(n11182), .O(n9139) );
  ND3CHD U6765 ( .I1(n12596), .I2(n10369), .I3(n10837), .O(n10382) );
  NR2EHD U6766 ( .I1(n12922), .I2(n12921), .O(n12925) );
  ND2DHD U6767 ( .I1(n8920), .I2(n6643), .O(n12883) );
  NR2CHD U6768 ( .I1(n8716), .I2(n13587), .O(n8752) );
  NR2CHD U6769 ( .I1(n9048), .I2(n11283), .O(n11289) );
  NR2GHD U6770 ( .I1(n10236), .I2(n12342), .O(n10235) );
  ND2CHD U6771 ( .I1(n7022), .I2(n7751), .O(n10826) );
  NR2GHD U6772 ( .I1(n9124), .I2(n9973), .O(n9123) );
  NR2CHD U6773 ( .I1(n10805), .I2(n7322), .O(n6994) );
  NR2EHD U6774 ( .I1(n11532), .I2(n8094), .O(n8093) );
  NR2GHD U6775 ( .I1(n10357), .I2(n10356), .O(n9457) );
  NR2CHD U6776 ( .I1(n13388), .I2(n9246), .O(n9245) );
  NR2GHD U6777 ( .I1(n7554), .I2(n7553), .O(n7867) );
  NR2CHD U6778 ( .I1(n12353), .I2(n12417), .O(n9281) );
  ND2DHD U6779 ( .I1(n9104), .I2(n7305), .O(n11384) );
  INVDHD U6780 ( .I(n11057), .O(n9535) );
  NR2CHD U6781 ( .I1(n8453), .I2(n6945), .O(n7373) );
  INVGHD U6782 ( .I(n10177), .O(n6891) );
  ND2DHD U6783 ( .I1(n11028), .I2(n12741), .O(n8456) );
  ND2CHD U6784 ( .I1(n11413), .I2(n8330), .O(n8481) );
  NR2BHD U6785 ( .I1(n12386), .I2(n12385), .O(n12387) );
  NR2GHD U6786 ( .I1(n11650), .I2(n8340), .O(n14078) );
  ND2CHD U6787 ( .I1(n8221), .I2(n11750), .O(n11754) );
  ND2DHD U6788 ( .I1(n13491), .I2(n8248), .O(n10194) );
  NR2BHD U6789 ( .I1(n11224), .I2(n11223), .O(n9583) );
  NR2CHD U6790 ( .I1(n8570), .I2(n10886), .O(n8569) );
  INVDHD U6791 ( .I(n11264), .O(n10015) );
  ND2CHD U6792 ( .I1(n7745), .I2(n6967), .O(n10819) );
  NR2EHD U6793 ( .I1(n11551), .I2(n11159), .O(n11534) );
  ND2HHD U6794 ( .I1(n13482), .I2(n9490), .O(n9487) );
  NR2BHD U6795 ( .I1(n12169), .I2(n12170), .O(n12177) );
  INVGHD U6796 ( .I(n7899), .O(n10989) );
  NR2GHD U6797 ( .I1(n12429), .I2(n12428), .O(n12430) );
  INVDHD U6798 ( .I(n6718), .O(n6695) );
  NR2EHD U6799 ( .I1(n13435), .I2(n12440), .O(n9722) );
  INVCKGHD U6800 ( .I(n12763), .O(n6783) );
  NR2EHD U6801 ( .I1(n11847), .I2(n7501), .O(n11851) );
  NR2CHD U6802 ( .I1(n11031), .I2(n10177), .O(n11032) );
  ND3CHD U6803 ( .I1(n11206), .I2(n11216), .I3(n9663), .O(n11207) );
  NR2BHD U6804 ( .I1(n8843), .I2(n11731), .O(n8838) );
  ND2DHD U6805 ( .I1(n13596), .I2(n12920), .O(n7553) );
  BUFJHD U6806 ( .I(n6820), .O(n7109) );
  INVGHD U6807 ( .I(n13828), .O(n7019) );
  AN2EHD U6808 ( .I1(n11553), .I2(n11155), .O(n11272) );
  AN2EHD U6809 ( .I1(n9832), .I2(n13133), .O(n13135) );
  AN2EHD U6810 ( .I1(n10798), .I2(n7172), .O(n6992) );
  BUFIHD U6811 ( .I(n12479), .O(n6588) );
  AN2EHD U6812 ( .I1(n12192), .I2(n14082), .O(n11761) );
  ND2DHD U6813 ( .I1(n9639), .I2(n8866), .O(n7554) );
  ND2DHD U6814 ( .I1(n8235), .I2(n8208), .O(n12633) );
  NR2CHD U6815 ( .I1(n9036), .I2(n12724), .O(n8462) );
  ND2DHD U6816 ( .I1(n12181), .I2(n8253), .O(n11844) );
  ND2DHD U6817 ( .I1(n13643), .I2(n13550), .O(n8844) );
  BUFIHD U6818 ( .I(n13818), .O(n6684) );
  BUFJHD U6819 ( .I(n9443), .O(n6520) );
  ND2DHD U6820 ( .I1(n11531), .I2(n9627), .O(n12470) );
  ND3CHD U6821 ( .I1(n12306), .I2(n13810), .I3(n7440), .O(n8841) );
  AN2EHD U6822 ( .I1(n8018), .I2(n12766), .O(n8373) );
  ND2DHD U6823 ( .I1(n11292), .I2(n9298), .O(n11532) );
  ND2DHD U6824 ( .I1(n12468), .I2(n6894), .O(n11143) );
  BUFJHD U6825 ( .I(n11297), .O(n9031) );
  ND3CHD U6826 ( .I1(n13182), .I2(n7382), .I3(n13603), .O(n7959) );
  INVGHD U6827 ( .I(n12813), .O(n10283) );
  ND3CHD U6828 ( .I1(n9300), .I2(n9152), .I3(n13680), .O(n11789) );
  BUFCKHHD U6829 ( .I(n13114), .O(n9596) );
  INVCKGHD U6830 ( .I(n12359), .O(n11937) );
  INVGHD U6831 ( .I(n10240), .O(n10237) );
  ND3CHD U6832 ( .I1(n12498), .I2(n12497), .I3(n8179), .O(n12499) );
  INVIHD U6833 ( .I(n12398), .O(n12399) );
  BUFKHD U6834 ( .I(n7450), .O(n6682) );
  INVGHD U6835 ( .I(n11508), .O(n10177) );
  ND2CHD U6836 ( .I1(n12856), .I2(n12864), .O(n12793) );
  NR2CHD U6837 ( .I1(n12240), .I2(n12237), .O(n7565) );
  NR2GHD U6838 ( .I1(n6988), .I2(n10021), .O(n7183) );
  ND2HHD U6839 ( .I1(n13596), .I2(n13590), .O(n13584) );
  ND2CHD U6840 ( .I1(n10207), .I2(n7223), .O(n10821) );
  ND2DHD U6841 ( .I1(n9104), .I2(n12766), .O(n11487) );
  NR2BHD U6842 ( .I1(n10630), .I2(n10796), .O(n10369) );
  ND2CHD U6843 ( .I1(n12247), .I2(n12331), .O(n8673) );
  INVGHD U6844 ( .I(n11731), .O(n13819) );
  NR2GHD U6845 ( .I1(n12211), .I2(n9695), .O(n14079) );
  AN2CHD U6846 ( .I1(n7499), .I2(n10073), .O(n12771) );
  INVGHD U6847 ( .I(n12965), .O(n12235) );
  ND2DHD U6848 ( .I1(n11364), .I2(n11411), .O(n8869) );
  AN2CHD U6849 ( .I1(n13022), .I2(n12364), .O(n6984) );
  NR2EHD U6850 ( .I1(n7678), .I2(n7684), .O(n7683) );
  INVJHD U6851 ( .I(n6574), .O(n8350) );
  NR2EHD U6852 ( .I1(n7706), .I2(n11025), .O(n11029) );
  INVGHD U6853 ( .I(n7504), .O(n6619) );
  NR2EHD U6854 ( .I1(n12504), .I2(n9294), .O(n9293) );
  ND2DHD U6855 ( .I1(n11365), .I2(n11349), .O(n11495) );
  BUFIHD U6856 ( .I(n12427), .O(n8876) );
  NR2GHD U6857 ( .I1(n11635), .I2(n12187), .O(n11636) );
  OR3EHD U6858 ( .I1(n7024), .I2(n12624), .I3(n10265), .O(n10264) );
  ND3CHD U6859 ( .I1(n9505), .I2(n11617), .I3(n8190), .O(n11618) );
  INVKHD U6860 ( .I(n11300), .O(n11312) );
  NR2EHD U6861 ( .I1(n11436), .I2(n11435), .O(n11557) );
  NR2EHD U6862 ( .I1(n7695), .I2(n9217), .O(n7692) );
  ND3CHD U6863 ( .I1(n8194), .I2(n7033), .I3(n9521), .O(n10736) );
  NR2EHD U6864 ( .I1(n12504), .I2(n9231), .O(n11426) );
  ND3CHD U6865 ( .I1(n9311), .I2(n7393), .I3(n13421), .O(n13002) );
  ND3CHD U6866 ( .I1(n6653), .I2(n6651), .I3(n13022), .O(n12964) );
  ND2CHD U6867 ( .I1(n7309), .I2(n11485), .O(n10537) );
  ND2DHD U6868 ( .I1(n13076), .I2(n12208), .O(n11621) );
  INVGHD U6869 ( .I(n7728), .O(n12872) );
  NR2EHD U6870 ( .I1(n8593), .I2(n8978), .O(n8592) );
  ND2CHD U6871 ( .I1(n7580), .I2(n12611), .O(n11248) );
  NR2GHD U6872 ( .I1(n8823), .I2(n10572), .O(n9111) );
  INVGHD U6873 ( .I(n12928), .O(n10135) );
  INVDHD U6874 ( .I(n11737), .O(n11721) );
  ND2DHD U6875 ( .I1(n13084), .I2(n13083), .O(n13087) );
  ND2CHD U6876 ( .I1(n13471), .I2(n8190), .O(n8668) );
  NR2BHD U6877 ( .I1(n12052), .I2(n12272), .O(n10009) );
  ND2CHD U6878 ( .I1(n9119), .I2(n13459), .O(n13033) );
  INVHHD U6879 ( .I(n6697), .O(n8221) );
  NR2GHD U6880 ( .I1(n7026), .I2(n9296), .O(n12476) );
  ND3CHD U6881 ( .I1(n13025), .I2(n9632), .I3(n9846), .O(n13026) );
  ND2HHD U6882 ( .I1(n12451), .I2(n11192), .O(n7899) );
  INVCKGHD U6883 ( .I(n10535), .O(n10536) );
  ND2DHD U6884 ( .I1(n9176), .I2(n13833), .O(n13834) );
  ND2HHD U6885 ( .I1(n12598), .I2(n6987), .O(n12532) );
  BUFHHD U6886 ( .I(n12419), .O(n9026) );
  ND2DHD U6887 ( .I1(n8339), .I2(n7304), .O(n11549) );
  INVGHD U6888 ( .I(n7395), .O(n13212) );
  ND2CHD U6889 ( .I1(n6677), .I2(n11814), .O(n13808) );
  ND2HHD U6890 ( .I1(n10992), .I2(n10991), .O(n9388) );
  NR2BHD U6891 ( .I1(n7207), .I2(n10069), .O(n6922) );
  INVJHD U6892 ( .I(n12322), .O(n7124) );
  ND2HHD U6893 ( .I1(n9520), .I2(n7008), .O(n9728) );
  OR2HHD U6894 ( .I1(n12196), .I2(n7502), .O(n7501) );
  INVGHD U6895 ( .I(n13427), .O(n9246) );
  ND2CHD U6896 ( .I1(n12705), .I2(n12704), .O(n12706) );
  NR2CHD U6897 ( .I1(n10223), .I2(n10224), .O(n10222) );
  NR2CHD U6898 ( .I1(n10621), .I2(n10620), .O(n10622) );
  NR2CHD U6899 ( .I1(n9153), .I2(n10261), .O(n11718) );
  NR2GHD U6900 ( .I1(n9404), .I2(n12971), .O(n12972) );
  ND3CHD U6901 ( .I1(n8153), .I2(n9674), .I3(n12383), .O(n12265) );
  NR2CHD U6902 ( .I1(n13029), .I2(n12957), .O(n12958) );
  NR2CHD U6903 ( .I1(n11900), .I2(n11899), .O(n11901) );
  BUFEHD U6904 ( .I(n7967), .O(n7966) );
  INVDHD U6905 ( .I(n10899), .O(n8915) );
  INVGHD U6906 ( .I(n6570), .O(n13218) );
  INVDHD U6907 ( .I(n13811), .O(n8839) );
  AN2CHD U6908 ( .I1(n13372), .I2(n9342), .O(n9341) );
  ND3CHD U6909 ( .I1(n11522), .I2(n11155), .I3(n10990), .O(n11435) );
  BUFGHD U6910 ( .I(n12869), .O(n7155) );
  ND2DHD U6911 ( .I1(n11295), .I2(n11459), .O(n11424) );
  BUFCKIHD U6912 ( .I(n14051), .O(n6641) );
  BUFIHD U6913 ( .I(n12735), .O(n8463) );
  AN2EHD U6914 ( .I1(n7942), .I2(n12123), .O(n8135) );
  AN2CHD U6915 ( .I1(n13440), .I2(n13419), .O(n13025) );
  AN2CHD U6916 ( .I1(n8962), .I2(n8888), .O(n8546) );
  AN2EHD U6917 ( .I1(n13582), .I2(n13614), .O(n7010) );
  AN2EHD U6918 ( .I1(n9770), .I2(n12945), .O(n12027) );
  AN2EHD U6919 ( .I1(n10959), .I2(n12868), .O(n8545) );
  ND2DHD U6920 ( .I1(n8866), .I2(n13590), .O(n10223) );
  ND3CHD U6921 ( .I1(n12338), .I2(n13004), .I3(n9398), .O(n12413) );
  BUFIHD U6922 ( .I(n12553), .O(n9104) );
  NR2EHD U6923 ( .I1(n13029), .I2(n13030), .O(n9252) );
  ND3CHD U6924 ( .I1(n11553), .I2(n12469), .I3(n11155), .O(n10701) );
  ND2DHD U6925 ( .I1(n7539), .I2(n11368), .O(n7706) );
  INVDHD U6926 ( .I(n13222), .O(n7027) );
  INVKHD U6927 ( .I(n9695), .O(n7594) );
  ND2CHD U6928 ( .I1(n10828), .I2(n12858), .O(n12849) );
  INVHHD U6929 ( .I(n9152), .O(n10261) );
  BUFCKHHD U6930 ( .I(n7487), .O(n7486) );
  NR2EHD U6931 ( .I1(n8029), .I2(n11752), .O(n9316) );
  ND2CHD U6932 ( .I1(n12559), .I2(n12768), .O(n7207) );
  INVGHD U6933 ( .I(n12970), .O(n12971) );
  BUFKHD U6934 ( .I(n13628), .O(n6543) );
  OR2EHD U6935 ( .I1(n12856), .I2(n12864), .O(n12840) );
  ND2CHD U6936 ( .I1(n9012), .I2(n9116), .O(n11436) );
  ND2DHD U6937 ( .I1(n11506), .I2(n11333), .O(n11025) );
  BUFJHD U6938 ( .I(n13602), .O(n9463) );
  BUFHHD U6939 ( .I(n9612), .O(n6677) );
  INVCKLHD U6940 ( .I(n9446), .O(n11307) );
  INVKHD U6941 ( .I(n7870), .O(n13211) );
  BUFKHD U6942 ( .I(n12655), .O(n9663) );
  BUFCKIHD U6943 ( .I(n7657), .O(n6789) );
  ND2CHD U6944 ( .I1(n12383), .I2(n11995), .O(n12384) );
  NR2EHD U6945 ( .I1(n13216), .I2(n13241), .O(n8329) );
  ND2HHD U6946 ( .I1(n13510), .I2(n13838), .O(n13809) );
  ND2DHD U6947 ( .I1(n7118), .I2(n13099), .O(n8998) );
  NR2CHD U6948 ( .I1(n12966), .I2(n12967), .O(n12969) );
  INVKHD U6949 ( .I(n6518), .O(n11263) );
  ND2DHD U6950 ( .I1(n7365), .I2(n12619), .O(n7642) );
  NR2EHD U6951 ( .I1(n10450), .I2(n7457), .O(n7456) );
  NR2GHD U6952 ( .I1(n10021), .I2(n7182), .O(n9708) );
  INVKHD U6953 ( .I(n8175), .O(n12898) );
  INVMHD U6954 ( .I(n13097), .O(n13083) );
  AN2EHD U6955 ( .I1(n6894), .I2(n9218), .O(n8436) );
  INVJHD U6956 ( .I(n7177), .O(n7178) );
  AN2EHD U6957 ( .I1(n7307), .I2(n12752), .O(n12728) );
  AN2EHD U6958 ( .I1(n12312), .I2(n13805), .O(n13660) );
  ND2DHD U6959 ( .I1(n8223), .I2(n12383), .O(n12276) );
  INVKHD U6960 ( .I(n9086), .O(n11376) );
  AN2EHD U6961 ( .I1(n12309), .I2(n13642), .O(n12310) );
  INVGHD U6962 ( .I(n12454), .O(n7026) );
  ND2DHD U6963 ( .I1(n12930), .I2(n11995), .O(n13207) );
  AN2CHD U6964 ( .I1(n12726), .I2(n12737), .O(n8430) );
  AN2CHD U6965 ( .I1(n12163), .I2(n12296), .O(n8252) );
  ND2DHD U6966 ( .I1(n9608), .I2(n7032), .O(n12217) );
  AN2EHD U6967 ( .I1(n11546), .I2(n9443), .O(n11419) );
  NR2EHD U6968 ( .I1(n12359), .I2(n12360), .O(n12362) );
  AN2CHD U6969 ( .I1(n11459), .I2(n9034), .O(n8246) );
  NR2BHD U6970 ( .I1(n7675), .I2(n7039), .O(n11325) );
  NR2EHD U6971 ( .I1(n7469), .I2(n7468), .O(n7467) );
  NR2EHD U6972 ( .I1(n13423), .I2(n13375), .O(n12414) );
  AN2EHD U6973 ( .I1(n12999), .I2(n13365), .O(n13001) );
  AN2EHD U6974 ( .I1(n10961), .I2(n8232), .O(n8240) );
  ND3CHD U6975 ( .I1(n7835), .I2(n13821), .I3(n13804), .O(n8753) );
  AN2EHD U6976 ( .I1(n8193), .I2(n12677), .O(n6968) );
  ND2CHD U6977 ( .I1(n11417), .I2(n11274), .O(n10704) );
  AN2EHD U6978 ( .I1(n10073), .I2(n12742), .O(n10528) );
  INVGHD U6979 ( .I(n6673), .O(n6921) );
  INVJHD U6980 ( .I(n11260), .O(n8138) );
  NR2EHD U6981 ( .I1(n11075), .I2(n11076), .O(n11077) );
  OR2EHD U6982 ( .I1(n9385), .I2(n10763), .O(n8492) );
  NR2EHD U6983 ( .I1(n7246), .I2(n7882), .O(n7881) );
  BUFMHD U6984 ( .I(n13208), .O(n6529) );
  INVLHD U6985 ( .I(n11814), .O(n13836) );
  INVGHD U6986 ( .I(n9342), .O(n8884) );
  NR2EHD U6987 ( .I1(n13011), .I2(n13449), .O(n12354) );
  ND2DHD U6988 ( .I1(n12743), .I2(n7028), .O(n11398) );
  BUFJHD U6989 ( .I(n13401), .O(n9589) );
  OR3EHD U6990 ( .I1(n11156), .I2(n11157), .I3(n11158), .O(n11163) );
  NR2EHD U6991 ( .I1(n8650), .I2(n11619), .O(n7369) );
  NR2EHD U6992 ( .I1(n10784), .I2(n10870), .O(n10786) );
  BUFIHD U6993 ( .I(n13420), .O(n9632) );
  NR2GHD U6994 ( .I1(n12346), .I2(n10126), .O(n13367) );
  ND2DHD U6995 ( .I1(n6970), .I2(n10958), .O(n8968) );
  NR2GHD U6996 ( .I1(n13670), .I2(n12081), .O(n9199) );
  NR2EHD U6997 ( .I1(n9351), .I2(n12579), .O(n11407) );
  ND2DHD U6998 ( .I1(n11510), .I2(n12553), .O(n10516) );
  INVGHD U6999 ( .I(n11280), .O(n9019) );
  ND2DHD U7000 ( .I1(n7247), .I2(n12869), .O(n10886) );
  ND2DHD U7001 ( .I1(n13373), .I2(n9093), .O(n13006) );
  ND2CHD U7002 ( .I1(n12766), .I2(n7539), .O(n11045) );
  ND2CHD U7003 ( .I1(n12868), .I2(n8337), .O(n10816) );
  ND2CHD U7004 ( .I1(n8204), .I2(n13231), .O(n14062) );
  BUFJHD U7005 ( .I(n13572), .O(n7031) );
  INVJHD U7006 ( .I(n12425), .O(n12353) );
  INVGHD U7007 ( .I(n8029), .O(n11626) );
  ND2CHD U7008 ( .I1(n12419), .I2(n13021), .O(n11899) );
  NR2EHD U7009 ( .I1(n12666), .I2(n12665), .O(n8140) );
  INVDHD U7010 ( .I(n9119), .O(n9234) );
  ND2CHD U7011 ( .I1(n11079), .I2(n9191), .O(n11081) );
  INVHHD U7012 ( .I(n8016), .O(n7681) );
  INVGHD U7013 ( .I(n6605), .O(n11625) );
  INVGHD U7014 ( .I(n7963), .O(n6835) );
  BUFEHD U7015 ( .I(n6801), .O(n6570) );
  ND2DHD U7016 ( .I1(n7454), .I2(n8511), .O(n8969) );
  ND2DHD U7017 ( .I1(n7606), .I2(n11233), .O(n10856) );
  ND2DHD U7018 ( .I1(n12173), .I2(n8178), .O(n13538) );
  ND2HHD U7019 ( .I1(n7187), .I2(n11254), .O(n12540) );
  INVCKGHD U7020 ( .I(n11279), .O(n9229) );
  NR2CHD U7021 ( .I1(n8917), .I2(n10756), .O(n9963) );
  NR2GHD U7022 ( .I1(n12874), .I2(n7747), .O(n7746) );
  NR2GHD U7023 ( .I1(n9197), .I2(n10143), .O(n10142) );
  ND2HHD U7024 ( .I1(n12999), .I2(n12364), .O(n13422) );
  INVGHD U7025 ( .I(n7929), .O(n13806) );
  ND2CHD U7026 ( .I1(n9593), .I2(n10618), .O(n10621) );
  ND2CHD U7027 ( .I1(n10889), .I2(n8145), .O(n8144) );
  BUFHHD U7028 ( .I(n12880), .O(n10207) );
  INVDHD U7029 ( .I(n11403), .O(n11341) );
  ND2HHD U7030 ( .I1(n12622), .I2(n12617), .O(n10630) );
  BUFJHD U7031 ( .I(n9462), .O(n9230) );
  NR2EHD U7032 ( .I1(MODE_1), .I2(KEYSET), .O(n10909) );
  INVGHD U7033 ( .I(n7229), .O(n7522) );
  INVGHD U7034 ( .I(n14053), .O(n8878) );
  INVHHD U7035 ( .I(n13223), .O(n9920) );
  NR2CHD U7036 ( .I1(n12122), .I2(n10129), .O(n7408) );
  ND2HHD U7037 ( .I1(n7366), .I2(n8615), .O(n8909) );
  INVJHD U7038 ( .I(n9682), .O(n10483) );
  NR2EHD U7039 ( .I1(n12034), .I2(n12033), .O(n12038) );
  NR2BHD U7040 ( .I1(n8926), .I2(n10214), .O(n8925) );
  INVGHD U7041 ( .I(n6640), .O(n8442) );
  NR2EHD U7042 ( .I1(n7441), .I2(n12367), .O(n12368) );
  BUFGHD U7043 ( .I(n12656), .O(n7154) );
  BUFHHD U7044 ( .I(n13383), .O(n9548) );
  BUFLHD U7045 ( .I(n6817), .O(n9687) );
  INVJHD U7046 ( .I(n12747), .O(n12778) );
  BUFIHD U7047 ( .I(n11337), .O(n9607) );
  BUFMHD U7048 ( .I(n11019), .O(n8607) );
  BUFJHD U7049 ( .I(n13399), .O(n9587) );
  INVGHD U7050 ( .I(n10021), .O(n7184) );
  INVDHD U7051 ( .I(n14051), .O(n8650) );
  AN2CHD U7052 ( .I1(n7223), .I2(n9003), .O(n7222) );
  BUFLHD U7053 ( .I(n13005), .O(n7139) );
  INVDHD U7054 ( .I(n10849), .O(n10784) );
  INVDHD U7055 ( .I(n10907), .O(n8509) );
  ND2DHD U7056 ( .I1(n9811), .I2(n11812), .O(n13811) );
  INVCHD U7057 ( .I(n11948), .O(n13432) );
  INVJHD U7058 ( .I(n12640), .O(n7182) );
  ND2HHD U7059 ( .I1(n9581), .I2(n10760), .O(n12869) );
  ND2DHD U7060 ( .I1(n7954), .I2(n9886), .O(n7465) );
  ND2DHD U7061 ( .I1(n12453), .I2(n9012), .O(n9292) );
  ND2DHD U7062 ( .I1(n12935), .I2(n12280), .O(n7466) );
  AN2EHD U7063 ( .I1(n9084), .I2(n13447), .O(n12956) );
  AN2HHD U7064 ( .I1(n10095), .I2(n8185), .O(n13576) );
  INVGHD U7065 ( .I(n14082), .O(n11619) );
  BUFLHD U7066 ( .I(n11521), .O(n9034) );
  ND2DHD U7067 ( .I1(n10296), .I2(n13487), .O(n9489) );
  BUFCKIHD U7068 ( .I(n12713), .O(n6706) );
  BUFJHD U7069 ( .I(n11512), .O(n7152) );
  BUFCKIHD U7070 ( .I(n9759), .O(n6694) );
  ND2DHD U7071 ( .I1(n9809), .I2(n7254), .O(n9808) );
  ND2HHD U7072 ( .I1(n13401), .I2(n9398), .O(n13015) );
  ND2HHD U7073 ( .I1(n7292), .I2(n7335), .O(n8254) );
  ND2HHD U7074 ( .I1(n7038), .I2(n9449), .O(n13019) );
  ND2HHD U7075 ( .I1(n12742), .I2(n11340), .O(n11392) );
  INVCHD U7076 ( .I(n11159), .O(n9295) );
  INVLHD U7077 ( .I(n13416), .O(n13426) );
  ND2CHD U7078 ( .I1(n7038), .I2(n7037), .O(n12426) );
  INVCHD U7079 ( .I(n8508), .O(n10214) );
  INVDHD U7080 ( .I(n6688), .O(n6687) );
  ND2DHD U7081 ( .I1(n10763), .I2(n9844), .O(n8879) );
  INVGHD U7082 ( .I(n12327), .O(n12328) );
  INVCHD U7083 ( .I(n12991), .O(n7269) );
  INVJHD U7084 ( .I(n10141), .O(n9197) );
  AN2EHD U7085 ( .I1(n12726), .I2(n11506), .O(n6944) );
  AN2CHD U7086 ( .I1(n12578), .I2(n7539), .O(n11412) );
  ND2HHD U7087 ( .I1(n7185), .I2(n7172), .O(n12634) );
  BUFIHD U7088 ( .I(n13194), .O(n6505) );
  ND2HHD U7089 ( .I1(n12291), .I2(n12031), .O(n13595) );
  AN2EHD U7090 ( .I1(n11410), .I2(n11411), .O(n6953) );
  INVJHD U7091 ( .I(n6644), .O(n13822) );
  BUFCKHHD U7092 ( .I(n12688), .O(n6647) );
  NR2EHD U7093 ( .I1(n13232), .I2(n9892), .O(n11758) );
  ND3CHD U7094 ( .I1(n9049), .I2(n7674), .I3(n7567), .O(n12754) );
  INVDHD U7095 ( .I(n12717), .O(n7457) );
  INVCHD U7096 ( .I(n11168), .O(n9297) );
  INVDHD U7097 ( .I(n9937), .O(n12950) );
  AN2EHD U7098 ( .I1(n12737), .I2(n11096), .O(n11097) );
  ND2HHD U7099 ( .I1(n7393), .I2(n12366), .O(n13449) );
  ND2HHD U7100 ( .I1(n12424), .I2(n7830), .O(n13400) );
  INVGHD U7101 ( .I(n13383), .O(n10126) );
  INVGHD U7102 ( .I(n13076), .O(n11630) );
  INVJHD U7103 ( .I(n7732), .O(n8615) );
  AN2CHD U7104 ( .I1(n12880), .I2(n10958), .O(n6975) );
  AN2CHD U7105 ( .I1(n12833), .I2(n7247), .O(n12806) );
  INVGHD U7106 ( .I(n7967), .O(n9488) );
  ND2CHD U7107 ( .I1(n12011), .I2(_i_CLEFIA128_keyL _39), .O(n9476) );
  ND2DHD U7108 ( .I1(n13510), .I2(n13805), .O(n11792) );
  BUFIHD U7109 ( .I(n10719), .O(n8858) );
  INVGHD U7110 ( .I(n13373), .O(n9928) );
  ND2HHD U7111 ( .I1(n13143), .I2(n13134), .O(n12122) );
  INVGHD U7112 ( .I(n7268), .O(n7267) );
  ND2DHD U7113 ( .I1(n6930), .I2(n12424), .O(n12323) );
  INVCKGHD U7114 ( .I(n12152), .O(n11776) );
  INVKHD U7115 ( .I(n11852), .O(n13489) );
  BUFJHD U7116 ( .I(n10965), .O(n6734) );
  AN2HHD U7117 ( .I1(n8832), .I2(n12150), .O(n13818) );
  BUFKHD U7118 ( .I(n7375), .O(n7374) );
  BUFIHD U7119 ( .I(n12952), .O(n9726) );
  ND2HHD U7120 ( .I1(n10141), .I2(n12089), .O(n12081) );
  NR2CHD U7121 ( .I1(n9441), .I2(n7886), .O(n7885) );
  ND2HHD U7122 ( .I1(n12656), .I2(n10855), .O(n7345) );
  INVCHD U7123 ( .I(n8235), .O(n9004) );
  INVGHD U7124 ( .I(n11409), .O(n8474) );
  BUFHHD U7125 ( .I(n12766), .O(n7679) );
  NR2CHD U7126 ( .I1(n6765), .I2(n6723), .O(n6784) );
  ND2DHD U7127 ( .I1(n9730), .I2(n9532), .O(n9460) );
  ND2HHD U7128 ( .I1(n9800), .I2(n11176), .O(n11429) );
  ND2HHD U7129 ( .I1(n8204), .I2(n7335), .O(n13471) );
  BUFIHD U7130 ( .I(n12846), .O(n7052) );
  ND2DHD U7131 ( .I1(n10794), .I2(n10793), .O(n11069) );
  INVKHD U7132 ( .I(n11406), .O(n9894) );
  INVGHD U7133 ( .I(n13613), .O(n12042) );
  BUFIHD U7134 ( .I(n8232), .O(n6716) );
  INVCKLHD U7135 ( .I(n9690), .O(n12609) );
  INVJHD U7136 ( .I(n8204), .O(n11609) );
  BUFJHD U7137 ( .I(n13191), .O(n7165) );
  ND2HHD U7138 ( .I1(n12327), .I2(n7038), .O(n9239) );
  BUFCKHHD U7139 ( .I(n7217), .O(n6615) );
  INVCKLHD U7140 ( .I(n6540), .O(n11508) );
  ND2HHD U7141 ( .I1(n12423), .I2(n9430), .O(n13371) );
  INVJHD U7142 ( .I(n6892), .O(n6893) );
  INVGHD U7143 ( .I(n10803), .O(n7318) );
  INVJHD U7144 ( .I(n8210), .O(n11615) );
  BUFJHD U7145 ( .I(n9800), .O(n9582) );
  INVMHD U7146 ( .I(n6804), .O(n6806) );
  NR2EHD U7147 ( .I1(n10450), .I2(n7455), .O(n8923) );
  INVCKGHD U7148 ( .I(n9898), .O(n11026) );
  ND2HHD U7149 ( .I1(n10760), .I2(n8916), .O(n12858) );
  INVHHD U7150 ( .I(n13216), .O(n13233) );
  INVGHD U7151 ( .I(n9185), .O(n9892) );
  INVGHD U7152 ( .I(n9194), .O(n6723) );
  INVKHD U7153 ( .I(n10794), .O(n6839) );
  ND2DHD U7154 ( .I1(n9811), .I2(n8178), .O(n11709) );
  INVJHD U7155 ( .I(n9741), .O(n10026) );
  ND2DHD U7156 ( .I1(n8113), .I2(n8006), .O(n11801) );
  INVLHD U7157 ( .I(n7908), .O(n10296) );
  INVCKLHD U7158 ( .I(n11230), .O(n11245) );
  INVGHD U7159 ( .I(n8962), .O(n8686) );
  NR2EHD U7160 ( .I1(n7890), .I2(n9092), .O(n7887) );
  INVHHD U7161 ( .I(n13829), .O(n7023) );
  INVJHD U7162 ( .I(n9165), .O(n13182) );
  INVHHD U7163 ( .I(n7340), .O(n9524) );
  INVCKLHD U7164 ( .I(n12846), .O(n12856) );
  ND2DHD U7165 ( .I1(n10884), .I2(n7720), .O(n12857) );
  ND2CHD U7166 ( .I1(n9626), .I2(n11181), .O(n6631) );
  INVKHD U7167 ( .I(n7206), .O(n10069) );
  ND2HHD U7168 ( .I1(n8977), .I2(n10728), .O(n8964) );
  ND2HHD U7169 ( .I1(n8237), .I2(n10690), .O(n11142) );
  INVGHD U7170 ( .I(n10960), .O(n7886) );
  ND2CHD U7171 ( .I1(n8215), .I2(n12794), .O(n12795) );
  ND2HHD U7172 ( .I1(n7291), .I2(n7078), .O(n13251) );
  INVJHD U7173 ( .I(n12578), .O(n7029) );
  ND2DHD U7174 ( .I1(n8194), .I2(n10965), .O(n7891) );
  INVDHD U7175 ( .I(n7083), .O(n8014) );
  INVLHD U7176 ( .I(n12424), .O(n12214) );
  INVLHD U7177 ( .I(n9007), .O(n8791) );
  NR2EHD U7178 ( .I1(n9744), .I2(n9062), .O(n9061) );
  INVKHD U7179 ( .I(n8191), .O(n9992) );
  INVHHD U7180 ( .I(n8938), .O(n10429) );
  BUFJHD U7181 ( .I(n11416), .O(n9017) );
  BUFEHD U7182 ( .I(n12748), .O(n7083) );
  INVDHD U7183 ( .I(n9383), .O(n10436) );
  INVLHD U7184 ( .I(n9810), .O(n12145) );
  AN2EHD U7185 ( .I1(n12561), .I2(n9801), .O(n6864) );
  INVDHD U7186 ( .I(n10737), .O(n10969) );
  INVKHD U7187 ( .I(n8218), .O(n6883) );
  INVKHD U7188 ( .I(n10252), .O(n8768) );
  INVKHD U7189 ( .I(n8218), .O(n12517) );
  INVMHD U7190 ( .I(n7969), .O(n12127) );
  ND2HHD U7191 ( .I1(n9699), .I2(n12129), .O(n12287) );
  INVHHD U7192 ( .I(n8194), .O(n10936) );
  INVDHD U7193 ( .I(n7038), .O(n9929) );
  INVKHD U7194 ( .I(n8095), .O(n7621) );
  ND2HHD U7195 ( .I1(n12424), .I2(n12251), .O(n12952) );
  ND2HHD U7196 ( .I1(n11049), .I2(n8188), .O(n11117) );
  AN2EHD U7197 ( .I1(n9099), .I2(n7132), .O(n11336) );
  INVDHD U7198 ( .I(n10966), .O(n9092) );
  NR2EHD U7199 ( .I1(n10090), .I2(n10431), .O(n9348) );
  INVCHD U7200 ( .I(n9214), .O(n12422) );
  AN2EHD U7201 ( .I1(n9841), .I2(n7132), .O(n6895) );
  BUFIHD U7202 ( .I(n9450), .O(n6562) );
  INVCHD U7203 ( .I(n7216), .O(n9532) );
  ND2HHD U7204 ( .I1(n7292), .I2(n9183), .O(n12192) );
  INVCKGHD U7205 ( .I(n11893), .O(n7037) );
  XNR2EHD U7206 ( .I1(_i_CLEFIA128_CON_T_xi _13), .I2(DOUT_62), .O(n10343));
  NR2EHD U7207 ( .I1(n10090), .I2(n9744), .O(n7244) );
  INVMHD U7208 ( .I(n7330), .O(n6804) );
  INVMHD U7209 ( .I(n9007), .O(n9680) );
  NR2EHD U7210 ( .I1(n7102), .I2(n8315), .O(n10884) );
  INVGHD U7211 ( .I(n9003), .O(n7455) );
  INVJHD U7212 ( .I(n12241), .O(n8887) );
  ND2CHD U7213 ( .I1(n7723), .I2(n10741), .O(n7722) );
  INVGHD U7214 ( .I(n8990), .O(n7968) );
  INVDHD U7215 ( .I(n7641), .O(n6785) );
  INVDHD U7216 ( .I(n11713), .O(n8113) );
  INVKHD U7217 ( .I(n12335), .O(n12324) );
  NR2CHD U7218 ( .I1(n6840), .I2(n11647), .O(n11763) );
  BUFNHD U7219 ( .I(n7336), .O(n7335) );
  INVNHD U7220 ( .I(n9349), .O(n10318) );
  ND2KHD U7221 ( .I1(n7036), .I2(n11713), .O(n13829) );
  NR2EHD U7222 ( .I1(n10090), .I2(n8207), .O(n12794) );
  INVLHD U7223 ( .I(n8095), .O(n8767) );
  OR2B1EHD U7224 ( .I1(n7014), .B1(n11505), .O(n11094) );
  BUFEHD U7225 ( .I(n9848), .O(n9620) );
  INVLHD U7226 ( .I(n8192), .O(n8193) );
  NR2GHD U7227 ( .I1(n8916), .I2(n8938), .O(n9993) );
  BUFJHD U7228 ( .I(n12830), .O(n7597) );
  BUFIHD U7229 ( .I(n10695), .O(n6765) );
  INVMHD U7230 ( .I(n10644), .O(n9007) );
  INVMHD U7231 ( .I(n7497), .O(n8188) );
  INVMHD U7232 ( .I(n10291), .O(n13442) );
  INVMHD U7233 ( .I(n11593), .O(n11766) );
  INVMHD U7234 ( .I(n8799), .O(n9435) );
  INVDHD U7235 ( .I(n9559), .O(n10088) );
  BUFMHD U7236 ( .I(n8224), .O(n6629) );
  XOR2HHD U7237 ( .I1(n8404), .I2(n7387), .O(n12335) );
  INVCHD U7238 ( .I(n10938), .O(n8960) );
  NR2GHD U7239 ( .I1(n12962), .I2(n9458), .O(n12241) );
  NR2GHD U7240 ( .I1(n10090), .I2(n12876), .O(n8936) );
  INVDHD U7241 ( .I(n11682), .O(n9095) );
  INVMHD U7242 ( .I(n6527), .O(n8218) );
  BUFCKHHD U7243 ( .I(n8212), .O(n6578) );
  BUFKHD U7244 ( .I(n6881), .O(n9777) );
  BUFHHD U7245 ( .I(n8164), .O(n7058) );
  ND2DHD U7246 ( .I1(n6775), .I2(n6773), .O(n10341) );
  BUFCKEHD U7247 ( .I(n12029), .O(n6810) );
  BUFNHD U7248 ( .I(n9887), .O(n9699) );
  INVIHD U7249 ( .I(n10090), .O(n9062) );
  INVKHD U7250 ( .I(n7016), .O(n7216) );
  BUFEHD U7251 ( .I(n7361), .O(n7360) );
  INVJHD U7252 ( .I(n12796), .O(n8192) );
  ND2CHD U7253 ( .I1(n6843), .I2(n6774), .O(n6773) );
  INVKHD U7254 ( .I(n7674), .O(n6876) );
  INVJHD U7255 ( .I(n9549), .O(n9480) );
  BUFJHD U7256 ( .I(n10636), .O(n6901) );
  NR2GHD U7257 ( .I1(n11991), .I2(n9187), .O(n11992) );
  BUFKHD U7258 ( .I(n8230), .O(n8903) );
  INVJHD U7259 ( .I(n10191), .O(n7703) );
  INVIHD U7260 ( .I(n8784), .O(n12962) );
  INVKHD U7261 ( .I(n6528), .O(n8799) );
  INVNHD U7262 ( .I(n7230), .O(n7723) );
  MUX2CHD U7263 ( .A(n10391), .B(n10390), .S(_i_CLEFIA128_keyL _78), .O(n10396) );
  MUX2CHD U7264 ( .A(n10575), .B(n10574), .S(_i_CLEFIA128_keyL _86), .O(n10580) );
  NR2CHD U7265 ( .I1(n9472), .I2(n7103), .O(n9471) );
  NR2GHD U7266 ( .I1(n10209), .I2(n10107), .O(n8167) );
  NR2EHD U7267 ( .I1(n14754), .I2(n7103), .O(n11597) );
  INVLHD U7268 ( .I(n11996), .O(n6881) );
  INVLHD U7269 ( .I(n9333), .O(n9332) );
  BUFMHD U7270 ( .I(n10767), .O(n10090) );
  INVJHD U7271 ( .I(n10259), .O(n7397) );
  ND2CHD U7272 ( .I1(n8224), .I2(_i_CLEFIA128_keyK _95), .O(n10345) );
  INVKHD U7273 ( .I(n10972), .O(n7042) );
  INVDHD U7274 ( .I(_i_CLEFIA128_keyL _63), .O(n6748) );
  OA112HHD U7275 ( .C1(n9414), .C2(n10032), .A1(n9413), .B1(n10028), .O(n8789));
  BUFMHD U7276 ( .I(n7977), .O(n7897) );
  INVGHD U7277 ( .I(n10431), .O(n7904) );
  BUFIHD U7278 ( .I(n11021), .O(n9750) );
  INVJHD U7279 ( .I(n10695), .O(n7053) );
  INVJHD U7280 ( .I(n6740), .O(n8201) );
  AN2EHD U7281 ( .I1(n7388), .I2(n7063), .O(n6634) );
  INVJHD U7282 ( .I(n8186), .O(n8187) );
  BUFCKIHD U7283 ( .I(n10442), .O(n6879) );
  INVKHD U7284 ( .I(n10107), .O(n9848) );
  ND2HHD U7285 ( .I1(n11896), .I2(n11904), .O(n11928) );
  INVJHD U7286 ( .I(n6523), .O(n10452) );
  INVGHD U7287 ( .I(n10266), .O(n7778) );
  AN2EHD U7288 ( .I1(n10338), .I2(n6776), .O(n6774) );
  INVJHD U7289 ( .I(n7783), .O(n6721) );
  INVJHD U7290 ( .I(n9844), .O(n9526) );
  NR2CHD U7291 ( .I1(n13984), .I2(n7103), .O(n10577) );
  INVLHD U7292 ( .I(n11896), .O(n11930) );
  INVJHD U7293 ( .I(n10145), .O(n9333) );
  INVDHD U7294 ( .I(_i_CLEFIA128_keyL _30), .O(n6776) );
  INVMHD U7295 ( .I(n10225), .O(n11628) );
  INVGHD U7296 ( .I(n10205), .O(n8411) );
  BUFJHD U7297 ( .I(n10445), .O(n9744) );
  NR2GHD U7298 ( .I1(n8207), .I2(n7338), .O(n9579) );
  ND2HHD U7299 ( .I1(n8115), .I2(n11685), .O(n12075) );
  INVMHD U7300 ( .I(n9206), .O(n9207) );
  BUFLHD U7301 ( .I(n7721), .O(n7720) );
  ND2CHD U7302 ( .I1(n11923), .I2(n6843), .O(n11925) );
  OR2B1EHD U7303 ( .I1(_i_CLEFIA128_keyK _15), .B1(n10337), .O(n10402) );
  INVNHD U7304 ( .I(n8315), .O(n10219) );
  INVLHD U7305 ( .I(n8136), .O(n7766) );
  XNR2HHD U7306 ( .I1(n10460), .I2(n8741), .O(n8230) );
  INVJHD U7307 ( .I(n7014), .O(n7567) );
  INVCKGHD U7308 ( .I(n6832), .O(n10479) );
  INVMHD U7309 ( .I(n7383), .O(n11707) );
  INVMHD U7310 ( .I(n12001), .O(n12914) );
  XNR2HHD U7311 ( .I1(n6890), .I2(n8717), .O(n6831) );
  INVCHD U7312 ( .I(n8378), .O(n7640) );
  ND2HHD U7313 ( .I1(n8133), .I2(n10446), .O(n10445) );
  INVMHD U7314 ( .I(n7389), .O(n10337) );
  XOR2EHD U7315 ( .I1(_i_CLEFIA128_CON_T_x _2), .I2(DOUT_113), .O(n6890) );
  XOR2CHD U7316 ( .I1(_i_CLEFIA128_CON_T_x _10), .I2(DOUT_106), .O(n6885) );
  INVMHD U7317 ( .I(n8206), .O(n10431) );
  OA12EHD U7318 ( .B1(n10254), .B2(n10310), .A1(_i_CLEFIA128_state_reg _1), .O(n10255) );
  ND3CHD U7319 ( .I1(n9411), .I2(n10030), .I3(n7389), .O(n10028) );
  INVMHD U7320 ( .I(n7225), .O(n10446) );
  INVDHD U7321 ( .I(n11587), .O(n9482) );
  INVDHD U7322 ( .I(n10308), .O(n10012) );
  ND2DHD U7323 ( .I1(n6834), .I2(n8159), .O(n8157) );
  INVGHD U7324 ( .I(n11870), .O(n11874) );
  XOR2EHD U7325 ( .I1(_i_CLEFIA128_CON_T_xi _11), .I2(DOUT_124), .O(n11587));
  XOR2EHD U7326 ( .I1(_i_CLEFIA128_CON_T_x _12), .I2(DOUT_59), .O(n10308) );
  ND2CHD U7327 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(_i_CLEFIA128_keyL _28), .O(n10254) );
  AN2EHD U7328 ( .I1(n9268), .I2(n11864), .O(n8290) );
  ND2CHD U7329 ( .I1(n11981), .I2(n7389), .O(n7201) );
  NR2EHD U7330 ( .I1(n7857), .I2(n9411), .O(n9410) );
  INVCHD U7331 ( .I(n10560), .O(n9906) );
  ND2HHD U7332 ( .I1(n11588), .I2(n7389), .O(n7643) );
  ND3CHD U7333 ( .I1(n8498), .I2(n9421), .I3(n6796), .O(n8496) );
  ND2DHD U7334 ( .I1(n8374), .I2(n15413), .O(n8676) );
  INVDHD U7335 ( .I(n6834), .O(n11980) );
  INVDHD U7336 ( .I(n9277), .O(n9275) );
  INVDHD U7337 ( .I(n9996), .O(n7763) );
  INVCKGHD U7338 ( .I(n9278), .O(n9276) );
  XOR2EHD U7339 ( .I1(_i_CLEFIA128_CON_T_xi_2 ), .I2(DOUT_51), .O(n10549) );
  XNR2EHD U7340 ( .I1(_i_CLEFIA128_CON_T_x _2), .I2(DOUT_49), .O(n8772) );
  XNR2CHD U7341 ( .I1(_i_CLEFIA128_CON_T_x _9), .I2(DOUT_32), .O(n6877) );
  XNR2CHD U7342 ( .I1(_i_CLEFIA128_CON_T_x _1), .I2(DOUT_48), .O(n10551) );
  XNR2CHD U7343 ( .I1(_i_CLEFIA128_CON_T_x _1), .I2(DOUT_40), .O(n10409) );
  INVDHD U7344 ( .I(_i_CLEFIA128_state_reg _1), .O(n9270) );
  XOR2CHD U7345 ( .I1(_i_CLEFIA128_CON_T_x _2), .I2(DOUT_41), .O(n8948) );
  NR2EHD U7346 ( .I1(n9721), .I2(n9168), .O(n9167) );
  ND2CHD U7347 ( .I1(n6622), .I2(_i_CLEFIA128_keyK _40), .O(n11865) );
  ND2CHD U7348 ( .I1(n8798), .I2(_i_CLEFIA128_keyL _69), .O(n9792) );
  ND2CHD U7349 ( .I1(n8798), .I2(_i_CLEFIA128_keyL _116), .O(n9394) );
  ND2DHD U7350 ( .I1(n8798), .I2(_i_CLEFIA128_keyL _107), .O(n11859) );
  ND2DHD U7351 ( .I1(n8798), .I2(_i_CLEFIA128_keyL _99), .O(n11967) );
  INVJHD U7352 ( .I(_i_CLEFIA128_keyL _52), .O(n15306) );
  INVGHD U7353 ( .I(_i_CLEFIA128_keyL _42), .O(n15413) );
  INVCHD U7354 ( .I(n10233), .O(n9949) );
  ND3CHD U7355 ( .I1(n11669), .I2(_i_CLEFIA128_rndcnt_reg _0), .I3(n15150), .O(n7541) );
  INVIHD U7356 ( .I(n6583), .O(n8319) );
  ND2HHD U7357 ( .I1(n8653), .I2(n6851), .O(n7414) );
  NR2GHD U7358 ( .I1(n8975), .I2(n7451), .O(n8940) );
  ND3CHD U7359 ( .I1(n8589), .I2(n11668), .I3(n8662), .O(n8661) );
  INVJHD U7360 ( .I(n6508), .O(n9395) );
  ND2DHD U7361 ( .I1(n8170), .I2(n11861), .O(n7560) );
  INVCHD U7362 ( .I(n9771), .O(n7434) );
  NR2EHD U7363 ( .I1(n8125), .I2(n8124), .O(n8123) );
  OA12EHD U7364 ( .B1(n8982), .B2(_i_CLEFIA128_keyK _101), .A1(n14405), .O(n11972) );
  INVLHD U7365 ( .I(_i_CLEFIA128_keyL _59), .O(n15078) );
  XOR2EHD U7366 ( .I1(_i_CLEFIA128_CON_T_x _10), .I2(DOUT_57), .O(n10233) );
  AN2EHD U7367 ( .I1(_i_CLEFIA128_keyK _36), .I2(_i_CLEFIA128_keyL _36), .O(n11963) );
  ND2CHD U7368 ( .I1(_i_CLEFIA128_keyK _27), .I2(_i_CLEFIA128_keyL _27), .O(n10306) );
  INVJHD U7369 ( .I(_i_CLEFIA128_keyL _34), .O(n15243) );
  ND3CHD U7370 ( .I1(n11977), .I2(_i_CLEFIA128_rndcnt_reg _0), .I3(n15280), .O(n7203) );
  NR2EHD U7371 ( .I1(n11888), .I2(n6899), .O(n10167) );
  ND2CHD U7372 ( .I1(_i_CLEFIA128_keyK _19), .I2(_i_CLEFIA128_keyL _19), .O(n10544) );
  ND2HHD U7373 ( .I1(n8039), .I2(_i_CLEFIA128_keyK _100), .O(n11964) );
  ND2CHD U7374 ( .I1(n9498), .I2(_i_CLEFIA128_keyL _125), .O(n9497) );
  XNR2HHD U7375 ( .I1(n8974), .I2(n10408), .O(n8973) );
  ND2CHD U7376 ( .I1(n8735), .I2(_i_CLEFIA128_rndcnt_reg _0), .O(n7780) );
  INVIHD U7377 ( .I(n9173), .O(n6796) );
  ND2DHD U7378 ( .I1(n8406), .I2(n10115), .O(n9203) );
  ND2DHD U7379 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(_i_CLEFIA128_keyK _49), .O(n8659) );
  INVDHD U7380 ( .I(n8944), .O(n8688) );
  INVLHD U7381 ( .I(_i_CLEFIA128_keyL _125), .O(n9502) );
  ND3CHD U7382 ( .I1(n8039), .I2(n15408), .I3(_i_CLEFIA128_keyK _64), .O(n8109) );
  XOR2EHD U7383 ( .I1(_i_CLEFIA128_CON_T_reg_4 ), .I2(DOUT_44), .O(n10411));
  ND3CHD U7384 ( .I1(n8797), .I2(n8902), .I3(_i_CLEFIA128_keyK _80), .O(n9201) );
  OR2HHD U7385 ( .I1(n7219), .I2(n9130), .O(n7006) );
  INVGHD U7386 ( .I(n14405), .O(n8691) );
  ND2DHD U7387 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(_i_CLEFIA128_keyL _44), .O(n11861) );
  ND2CHD U7388 ( .I1(_i_CLEFIA128_keyK _21), .I2(_i_CLEFIA128_keyL _21), .O(n10557) );
  ND2CHD U7389 ( .I1(_i_CLEFIA128_keyK _56), .I2(_i_CLEFIA128_keyL _56), .O(n11590) );
  ND2DHD U7390 ( .I1(_i_CLEFIA128_keyL _24), .I2(_i_CLEFIA128_keyK _24), .O(n7224) );
  ND2CHD U7391 ( .I1(n8798), .I2(_i_CLEFIA128_keyL _73), .O(n8946) );
  ND2CHD U7392 ( .I1(n8798), .I2(_i_CLEFIA128_keyL _67), .O(n10454) );
  ND2DHD U7393 ( .I1(_i_CLEFIA128_keyK _33), .I2(_i_CLEFIA128_keyL _33), .O(n11978) );
  ND2DHD U7394 ( .I1(_i_CLEFIA128_keyK _2), .I2(_i_CLEFIA128_keyL _2), .O(n10468) );
  ND2CHD U7395 ( .I1(n13778), .I2(_i_CLEFIA128_keyL _80), .O(n9200) );
  ND2HHD U7396 ( .I1(n8797), .I2(_i_CLEFIA128_keyK _113), .O(n11668) );
  INVJHD U7397 ( .I(_i_CLEFIA128_keyL _27), .O(n15247) );
  INVCKGHD U7398 ( .I(n10114), .O(n10115) );
  NR2EHD U7399 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(n9527), .O(n8947) );
  INVDHD U7400 ( .I(_i_CLEFIA128_keyL _61), .O(n6579) );
  ND2DHD U7401 ( .I1(n8797), .I2(_i_CLEFIA128_keyK _2), .O(n10466) );
  ND2CHD U7402 ( .I1(_i_CLEFIA128_keyK _58), .I2(_i_CLEFIA128_keyL _58), .O(n11572) );
  INVJHD U7403 ( .I(_i_CLEFIA128_keyL _50), .O(n15179) );
  INVJHD U7404 ( .I(_i_CLEFIA128_keyL _45), .O(n15073) );
  INVDHD U7405 ( .I(n10118), .O(n8574) );
  INVJHD U7406 ( .I(_i_CLEFIA128_keyL _53), .O(n14927) );
  ND2CHD U7407 ( .I1(n6745), .I2(_i_CLEFIA128_keyK _21), .O(n6744) );
  ND2HHD U7408 ( .I1(n8551), .I2(_i_CLEFIA128_state_reg _1), .O(n8559) );
  INVJHD U7409 ( .I(_i_CLEFIA128_keyL _57), .O(n15198) );
  INVJHD U7410 ( .I(_i_CLEFIA128_keyL _56), .O(n15140) );
  NR2GHD U7411 ( .I1(n6822), .I2(n8616), .O(n8928) );
  INVJHD U7412 ( .I(_i_CLEFIA128_keyL _20), .O(n15244) );
  INVGHD U7413 ( .I(_i_CLEFIA128_keyL _84), .O(n9130) );
  INVJHD U7414 ( .I(_i_CLEFIA128_keyL _24), .O(n14556) );
  ND2CHD U7415 ( .I1(n8039), .I2(_i_CLEFIA128_keyK _58), .O(n11570) );
  ND2DHD U7416 ( .I1(n8797), .I2(_i_CLEFIA128_keyK _4), .O(n10456) );
  INVKHD U7417 ( .I(_i_CLEFIA128_keyL _10), .O(n14991) );
  INVJHD U7418 ( .I(_i_CLEFIA128_keyL _51), .O(n15014) );
  INVJHD U7419 ( .I(_i_CLEFIA128_keyL _25), .O(n14953) );
  INVGHD U7420 ( .I(n6828), .O(n6829) );
  INVNHD U7421 ( .I(_i_CLEFIA128_keyL _3), .O(n15300) );
  INVJHD U7422 ( .I(_i_CLEFIA128_keyL _29), .O(n15176) );
  ND2DHD U7423 ( .I1(n6709), .I2(_i_CLEFIA128_keyK _12), .O(n6708) );
  INVJHD U7424 ( .I(_i_CLEFIA128_keyL _13), .O(n15242) );
  INVLHD U7425 ( .I(n14405), .O(n6850) );
  ND2KHD U7426 ( .I1(n15235), .I2(n15218), .O(n15228) );
  ND2KHD U7427 ( .I1(n15171), .I2(n15154), .O(n15164) );
  INVMHD U7428 ( .I(n8519), .O(n8521) );
  INVDHD U7429 ( .I(n8179), .O(n6750) );
  NR2IHD U7430 ( .I1(n7343), .I2(n8849), .O(n7974) );
  INVNHD U7431 ( .I(n8760), .O(n11834) );
  ND3EHD U7432 ( .I1(n9556), .I2(n13234), .I3(n13233), .O(n13236) );
  NR2GHD U7433 ( .I1(n10428), .I2(n7338), .O(n8961) );
  NR2GHD U7434 ( .I1(n8863), .I2(n8783), .O(n12763) );
  NR2EHD U7435 ( .I1(n12574), .I2(n11381), .O(n11386) );
  ND2DHD U7436 ( .I1(n14999), .I2(n7190), .O(n6199) );
  ND3CHD U7437 ( .I1(n14174), .I2(n14175), .I3(n14173), .O(n6211) );
  ND3CHD U7438 ( .I1(n7364), .I2(n9457), .I3(n10653), .O(n10654) );
  OR2B1CHD U7439 ( .I1(n11087), .B1(n10847), .O(n10676) );
  ND2HHD U7440 ( .I1(n8039), .I2(_i_CLEFIA128_keyK _27), .O(n7855) );
  AO12EHD U7441 ( .B1(n15200), .B2(n7043), .A1(n15199), .O(n6347) );
  NR2GHD U7442 ( .I1(n10710), .I2(n10727), .O(n9936) );
  OAI112BHD U7443 ( .C1(n6765), .C2(n9541), .A1(n11459), .B1(n12448), .O(n10697) );
  AN3HHD U7444 ( .I1(n9053), .I2(n11440), .I3(n6520), .O(n6999) );
  NR2EHD U7445 ( .I1(n13247), .I2(n13095), .O(n6771) );
  XNR2HHD U7446 ( .I1(n14169), .I2(n6808), .O(n8764) );
  XNR3EHD U7447 ( .I1(DOUT_8), .I2(n6889), .I3(n7110), .O(n7876) );
  XNR3EHD U7448 ( .I1(n10075), .I2(n7110), .I3(n13741), .O(n13742) );
  XNR2EHD U7449 ( .I1(n7110), .I2(n8774), .O(n9543) );
  INVGHD U7450 ( .I(n9434), .O(n9433) );
  NR2GHD U7451 ( .I1(n8849), .I2(n8355), .O(n7979) );
  XOR2HHD U7452 ( .I1(n8910), .I2(n7472), .O(n7471) );
  ND2DHD U7453 ( .I1(n15440), .I2(n11130), .O(n15430) );
  ND2DHD U7454 ( .I1(n15440), .I2(n15500), .O(n15444) );
  ND2HHD U7455 ( .I1(n7829), .I2(n7828), .O(n10172) );
  XOR2HHD U7456 ( .I1(n7955), .I2(n9409), .O(n14091) );
  ND2DHD U7457 ( .I1(n15193), .I2(n15500), .O(n13862) );
  OA12EHD U7458 ( .B1(n7191), .B2(n11129), .A1(n14998), .O(n7190) );
  ND2DHD U7459 ( .I1(n11948), .I2(n8229), .O(n10122) );
  XNR3EHD U7460 ( .I1(n9408), .I2(n14351), .I3(n8787), .O(n9407) );
  OR2EHD U7461 ( .I1(n15512), .I2(n15374), .O(n15370) );
  OR3EHD U7462 ( .I1(n13632), .I2(n13633), .I3(n13631), .O(n13637) );
  ND2DHD U7463 ( .I1(n15178), .I2(n11130), .O(n13567) );
  ND2DHD U7464 ( .I1(n8603), .I2(n8601), .O(n6205) );
  ND2HHD U7465 ( .I1(n10416), .I2(n10201), .O(n10200) );
  OAI12CHD U7466 ( .B1(n9895), .B2(n15416), .A1(n14663), .O(n6266) );
  ND2DHD U7467 ( .I1(n7616), .I2(n14836), .O(n6281) );
  AOI12HHD U7468 ( .B1(n15269), .B2(n15500), .A1(n14960), .O(n8354) );
  AOI12HHD U7469 ( .B1(n15269), .B2(n11130), .A1(n13163), .O(n7005) );
  OAI12CHD U7470 ( .B1(n15439), .B2(n15416), .A1(n14545), .O(n6325) );
  ND2HHD U7471 ( .I1(n13712), .I2(n13711), .O(n6103) );
  MUX2HHD U7472 ( .A(n13704), .B(n13703), .S(n14615), .O(n13712) );
  XNR2EHD U7473 ( .I1(n9816), .I2(n6852), .O(n10139) );
  INVLHD U7474 ( .I(n10188), .O(n10187) );
  BUFMHD U7475 ( .I(n14766), .O(n9089) );
  ND2HHD U7476 ( .I1(n9867), .I2(n7043), .O(n9866) );
  NR2CHD U7477 ( .I1(n11039), .I2(n11043), .O(n7263) );
  NR2EHD U7478 ( .I1(n7258), .I2(n7259), .O(n7257) );
  XNR2HHD U7479 ( .I1(n7213), .I2(n14995), .O(n7212) );
  ND2DHD U7480 ( .I1(n14813), .I2(n11130), .O(n13504) );
  INVMHD U7481 ( .I(n7680), .O(n11119) );
  INVKHD U7482 ( .I(n9737), .O(n10268) );
  ND2DHD U7483 ( .I1(n8007), .I2(n14841), .O(n6337) );
  ND2HHD U7484 ( .I1(n15520), .I2(n15506), .O(n15518) );
  NR2CHD U7485 ( .I1(n10689), .I2(n10688), .O(n10692) );
  NR2IHD U7486 ( .I1(n13610), .I2(n13611), .O(n13641) );
  ND2DHD U7487 ( .I1(n8307), .I2(n10044), .O(n6275) );
  XOR2HHD U7488 ( .I1(n14170), .I2(n10018), .O(n14013) );
  AO22CHD U7489 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _123), .B1(n15504), .B2(_i_CLEFIA128_keyK _59), .O(n8298) );
  ND3CHD U7490 ( .I1(n15448), .I2(n9149), .I3(n15447), .O(n6172) );
  ND2DHD U7491 ( .I1(n9151), .I2(n15500), .O(n9149) );
  ND2HHD U7492 ( .I1(n9151), .I2(n8263), .O(n9148) );
  ND2DHD U7493 ( .I1(n9151), .I2(n11130), .O(n9150) );
  NR2CHD U7494 ( .I1(n9944), .I2(n13813), .O(n13815) );
  ND2HHD U7495 ( .I1(n12267), .I2(n13122), .O(n7963) );
  XNR2KHD U7496 ( .I1(n6725), .I2(n7876), .O(n15392) );
  BUFMHD U7497 ( .I(n7985), .O(n6725) );
  XNR2KHD U7498 ( .I1(n14091), .I2(n7120), .O(n15193) );
  ND2HHD U7499 ( .I1(n15095), .I2(n8273), .O(n9714) );
  AN3HHD U7500 ( .I1(n9770), .I2(n13572), .I3(n12934), .O(n8324) );
  NR2IHD U7501 ( .I1(n7670), .I2(n8621), .O(n7669) );
  INVDHD U7502 ( .I(n13684), .O(n8621) );
  ND2HHD U7503 ( .I1(n7952), .I2(n15500), .O(n9999) );
  NR2GHD U7504 ( .I1(n10468), .I2(n6899), .O(n9787) );
  NR2EHD U7505 ( .I1(n12104), .I2(n12103), .O(n12105) );
  OA12EHD U7506 ( .B1(n7992), .B2(n8816), .A1(n8294), .O(n7295) );
  AN2HHD U7507 ( .I1(n8628), .I2(n7537), .O(n8803) );
  ND3CHD U7508 ( .I1(n9639), .I2(n13121), .I3(n13122), .O(n13123) );
  ND2HHD U7509 ( .I1(n9558), .I2(n13107), .O(n8790) );
  NR2GHD U7510 ( .I1(n13615), .I2(n13116), .O(n13119) );
  BUFNHD U7511 ( .I(n13591), .O(n9603) );
  XOR2HHD U7512 ( .I1(n13715), .I2(DOUT_1), .O(n13716) );
  BUFKHD U7513 ( .I(n14647), .O(n7082) );
  INVMHD U7514 ( .I(n7856), .O(n7866) );
  INVGHD U7515 ( .I(n10869), .O(n7151) );
  NR2EHD U7516 ( .I1(n8691), .I2(n11989), .O(n8690) );
  AN3B1EHD U7517 ( .I1(n14931), .I2(_i_CLEFIA128_keyK _68), .B1(n8798), .O(n7478) );
  NR2GHD U7518 ( .I1(n8798), .I2(n15058), .O(n7646) );
  ND2KHD U7519 ( .I1(n6504), .I2(n10185), .O(n9209) );
  ND2HHD U7520 ( .I1(n7914), .I2(n7915), .O(n6504) );
  NR2IHD U7521 ( .I1(n13158), .I2(n13159), .O(n13160) );
  OA12HHD U7522 ( .B1(n12130), .B2(n8990), .A1(n7417), .O(n12131) );
  INVKHD U7523 ( .I(n8155), .O(n12264) );
  ND2KHD U7524 ( .I1(n7433), .I2(n8396), .O(n7313) );
  ND2DHD U7525 ( .I1(n12637), .I2(n11079), .O(n10772) );
  NR2EHD U7526 ( .I1(n11249), .I2(n11248), .O(n11252) );
  NR2GHD U7527 ( .I1(n6813), .I2(n12544), .O(n12547) );
  ND3EHD U7528 ( .I1(n12477), .I2(n10987), .I3(n10986), .O(n11545) );
  AN2HHD U7529 ( .I1(n6998), .I2(n10119), .O(n12477) );
  NR2GHD U7530 ( .I1(n11716), .I2(n11717), .O(n11719) );
  AN2HHD U7531 ( .I1(n6506), .I2(n9732), .O(n13161) );
  OAI12CHD U7532 ( .B1(n6606), .B2(n13157), .A1(n6507), .O(n6506) );
  ND2HHD U7533 ( .I1(n9396), .I2(n14405), .O(n6508) );
  ND2KHD U7534 ( .I1(n6820), .I2(n6727), .O(n11395) );
  ND2HHD U7535 ( .I1(n6509), .I2(n8294), .O(n7429) );
  ND3EHD U7536 ( .I1(n8802), .I2(n7431), .I3(n6920), .O(n6509) );
  ND2KHD U7537 ( .I1(n12726), .I2(n12769), .O(n12757) );
  ND2HHD U7538 ( .I1(n7398), .I2(n7301), .O(n12769) );
  NR2CHD U7539 ( .I1(n7344), .I2(n9331), .O(n10879) );
  INVMHD U7540 ( .I(n10324), .O(n8854) );
  INVGHD U7541 ( .I(n11782), .O(n11723) );
  INVNHD U7542 ( .I(n6818), .O(n6819) );
  INVGHD U7543 ( .I(n6510), .O(n8251) );
  ND2HHD U7544 ( .I1(n8444), .I2(n7579), .O(n6510) );
  XOR2HHD U7545 ( .I1(_i_CLEFIA128_CON_T_x _10), .I2(DOUT_33), .O(n10464) );
  OR3HHD U7546 ( .I1(n6511), .I2(n7099), .I3(n8537), .O(n8535) );
  NR2GHD U7547 ( .I1(n6876), .I2(n11335), .O(n6511) );
  XOR2HHD U7548 ( .I1(n6874), .I2(n6815), .O(n10217) );
  ND3EHD U7549 ( .I1(n7514), .I2(n7512), .I3(n7509), .O(n6815) );
  ND2KHD U7550 ( .I1(n13121), .I2(n9998), .O(n9015) );
  ND2KHD U7551 ( .I1(n7968), .I2(n8183), .O(n13121) );
  ND3EHD U7552 ( .I1(n13829), .I2(n6512), .I3(n13820), .O(n12144) );
  INVGHD U7553 ( .I(n6513), .O(n6512) );
  ND2HHD U7554 ( .I1(n7537), .I2(n13643), .O(n6513) );
  ND2HHD U7555 ( .I1(n13037), .I2(n9311), .O(n6515) );
  INVGHD U7556 ( .I(n6516), .O(n6997) );
  ND2HHD U7557 ( .I1(n12620), .I2(n8235), .O(n6516) );
  AN2HHD U7558 ( .I1(n8916), .I2(n9348), .O(n8427) );
  INVGHD U7559 ( .I(n13051), .O(n12998) );
  INVQHD U7560 ( .I(n6517), .O(n12900) );
  INVNHD U7561 ( .I(n11993), .O(n6517) );
  INVCKLHD U7562 ( .I(n9774), .O(n7189) );
  AN2HHD U7563 ( .I1(_i_CLEFIA128_keyK _11), .I2(_i_CLEFIA128_keyL _11), .O(n8346) );
  INVIHD U7564 ( .I(n10827), .O(n6760) );
  ND3EHD U7565 ( .I1(n7514), .I2(n7509), .I3(n7512), .O(n6534) );
  ND2KHD U7566 ( .I1(n12640), .I2(n11079), .O(n6518) );
  NR2GHD U7567 ( .I1(n12300), .I2(n13662), .O(n12301) );
  MUX2HHD U7568 ( .A(n12817), .B(n12816), .S(n7998), .O(n12825) );
  BUFMHD U7569 ( .I(n11677), .O(n6872) );
  ND2KHD U7570 ( .I1(n6524), .I2(n11380), .O(n9036) );
  ND2KHD U7571 ( .I1(n8182), .I2(n12561), .O(n11380) );
  ND2HHD U7572 ( .I1(n6519), .I2(n13826), .O(n7050) );
  ND3EHD U7573 ( .I1(n7426), .I2(n7428), .I3(n6914), .O(n6519) );
  ND2KHD U7574 ( .I1(n8030), .I2(n10268), .O(n7170) );
  OR2KHD U7575 ( .I1(n10463), .I2(n6898), .O(n10245) );
  ND2KHD U7576 ( .I1(n7522), .I2(n8233), .O(n9553) );
  INVKHD U7577 ( .I(n6521), .O(n11415) );
  ND2HHD U7578 ( .I1(n7666), .I2(n7663), .O(n6521) );
  INVNHD U7579 ( .I(n9458), .O(n6909) );
  ND2KHD U7580 ( .I1(n8914), .I2(n10945), .O(n8919) );
  NR2IHD U7581 ( .I1(n8918), .I2(n8919), .O(n8489) );
  ND2HHD U7582 ( .I1(n6607), .I2(n13439), .O(n13012) );
  NR2IHD U7583 ( .I1(n13012), .I2(n13011), .O(n13013) );
  INVQHD U7584 ( .I(_i_CLEFIA128_keyL _106), .O(n8679) );
  ND3EHD U7585 ( .I1(n11876), .I2(n8589), .I3(n8679), .O(n8678) );
  ND3EHD U7586 ( .I1(n13005), .I2(n13373), .I3(n9084), .O(n9097) );
  INVKHD U7587 ( .I(n7970), .O(n6557) );
  XOR2HHD U7588 ( .I1(n8790), .I2(n8578), .O(n10004) );
  ND2HHD U7589 ( .I1(n10146), .I2(n12179), .O(n8578) );
  INVJHD U7590 ( .I(n10833), .O(n12516) );
  ND3EHD U7591 ( .I1(n8220), .I2(n11236), .I3(n7178), .O(n10833) );
  ND2KHD U7592 ( .I1(n7347), .I2(n6989), .O(n9331) );
  ND2KHD U7593 ( .I1(n8515), .I2(n12766), .O(n12738) );
  INVJHD U7594 ( .I(n6522), .O(n7585) );
  ND2KHD U7595 ( .I1(n7586), .I2(n7588), .O(n6522) );
  ND2HHD U7596 ( .I1(n8397), .I2(n7783), .O(n6523) );
  OA13EHD U7597 ( .B1(n7121), .B2(n8816), .B3(n12178), .A1(n13835), .O(n7293));
  ND3EHD U7598 ( .I1(n8341), .I2(n8579), .I3(n13833), .O(n8816) );
  ND2KHD U7599 ( .I1(n9041), .I2(n9547), .O(n14993) );
  INVJHD U7600 ( .I(n6681), .O(n7095) );
  NR2GHD U7601 ( .I1(n7731), .I2(n7729), .O(n7735) );
  ND2KHD U7602 ( .I1(n12517), .I2(n10318), .O(n12656) );
  ND2KHD U7603 ( .I1(n12651), .I2(n11253), .O(n9671) );
  ND2KHD U7604 ( .I1(n10318), .I2(n10874), .O(n11253) );
  ND2KHD U7605 ( .I1(n7398), .I2(n9694), .O(n6524) );
  ND3EHD U7606 ( .I1(n10051), .I2(n7383), .I3(n11679), .O(n6740) );
  NR2GHD U7607 ( .I1(n6525), .I2(n11854), .O(n9046) );
  OA13EHD U7608 ( .B1(n9445), .B2(n11846), .B3(n9354), .A1(n14087), .O(n6525));
  ND2KHD U7609 ( .I1(n12637), .I2(n12618), .O(n10848) );
  ND2KHD U7610 ( .I1(n9680), .I2(n10668), .O(n12637) );
  INVLHD U7611 ( .I(n11685), .O(n7777) );
  ND3EHD U7612 ( .I1(n6526), .I2(n10311), .I3(n10255), .O(n8874) );
  ND2HHD U7613 ( .I1(n10257), .I2(n6851), .O(n6526) );
  NR2EHD U7614 ( .I1(n10047), .I2(n12510), .O(n10046) );
  ND2KHD U7615 ( .I1(n12561), .I2(n8188), .O(n11333) );
  INVLHD U7616 ( .I(n9226), .O(n9923) );
  INVJHD U7617 ( .I(n10096), .O(n8875) );
  ND2KHD U7618 ( .I1(n10470), .I2(n6851), .O(n8525) );
  NR2IHD U7619 ( .I1(n8199), .I2(n12520), .O(n6527) );
  ND2KHD U7620 ( .I1(n10636), .I2(n7016), .O(n12520) );
  NR2GHD U7621 ( .I1(n11775), .I2(n7808), .O(n6528) );
  ND2KHD U7622 ( .I1(n7382), .I2(n12945), .O(n12107) );
  ND2KHD U7623 ( .I1(n8797), .I2(_i_CLEFIA128_keyK _115), .O(n11667) );
  NR2EHD U7624 ( .I1(n10946), .I2(n8532), .O(n8531) );
  NR2IHD U7625 ( .I1(n12113), .I2(n12112), .O(n12114) );
  NR2CHD U7626 ( .I1(n7895), .I2(n9507), .O(n9506) );
  ND3EHD U7627 ( .I1(n9523), .I2(n12856), .I3(n10825), .O(n9522) );
  NR2GHD U7628 ( .I1(n7941), .I2(n13662), .O(n7940) );
  ND3EHD U7629 ( .I1(n6530), .I2(n8072), .I3(n8069), .O(n11756) );
  INVCKGHD U7630 ( .I(n6531), .O(n6530) );
  ND2HHD U7631 ( .I1(n6737), .I2(n9646), .O(n6531) );
  ND3EHD U7632 ( .I1(n10493), .I2(n10494), .I3(_i_CLEFIA128_state_reg _1), .O(n10495) );
  AN3B1HHD U7633 ( .I1(n6589), .I2(n13222), .B1(n11844), .O(n11845) );
  OAI12CHD U7634 ( .B1(n10404), .B2(_i_CLEFIA128_keyL _15), .A1(n6532), .O(n10405) );
  OAI12CHD U7635 ( .B1(n7103), .B2(n14784), .A1(_i_CLEFIA128_keyL _15), .O(n6532) );
  NR2EHD U7636 ( .I1(n11330), .I2(n11331), .O(n11332) );
  ND2HHD U7637 ( .I1(n7109), .I2(n6952), .O(n10522) );
  INVMHD U7638 ( .I(n7410), .O(n11685) );
  ND3EHD U7639 ( .I1(n10241), .I2(n10240), .I3(n9019), .O(n9554) );
  NR2IHD U7640 ( .I1(n7894), .I2(n11556), .O(n10241) );
  INVJHD U7641 ( .I(n10619), .O(n6553) );
  INVJHD U7642 ( .I(n10619), .O(n11166) );
  XOR2HHD U7643 ( .I1(n6534), .I2(n9664), .O(n9818) );
  BUFMHD U7644 ( .I(n9772), .O(n6535) );
  INVGHD U7645 ( .I(n6536), .O(n8363) );
  ND2HHD U7646 ( .I1(n12899), .I2(n12290), .O(n6536) );
  ND3EHD U7647 ( .I1(n12401), .I2(n13183), .I3(n10080), .O(n12272) );
  ND2KHD U7648 ( .I1(n12291), .I2(n12129), .O(n13183) );
  BUFMHD U7649 ( .I(n9540), .O(n7952) );
  ND2KHD U7650 ( .I1(n12927), .I2(n13634), .O(n13111) );
  INVGHD U7651 ( .I(n6537), .O(n8098) );
  ND3EHD U7652 ( .I1(n8099), .I2(n14988), .I3(_i_CLEFIA128_rndcnt_reg _0), .O(n6537) );
  ND3EHD U7653 ( .I1(n12375), .I2(n9752), .I3(n6535), .O(n12380) );
  ND2HHD U7654 ( .I1(n9210), .I2(n9309), .O(n12147) );
  INVDHD U7655 ( .I(n9299), .O(n7918) );
  AN2HHD U7656 ( .I1(n10241), .I2(n7001), .O(n8413) );
  OA13EHD U7657 ( .B1(n8737), .B2(n12407), .B3(n13624), .A1(n13608), .O(n12408) );
  ND2HHD U7658 ( .I1(n12910), .I2(n9677), .O(n8737) );
  ND2HHD U7659 ( .I1(n13589), .I2(n12393), .O(n10133) );
  ND2HHD U7660 ( .I1(n12125), .I2(n11976), .O(n12393) );
  ND2KHD U7661 ( .I1(n8136), .I2(n10325), .O(n9774) );
  INVQHD U7662 ( .I(n6539), .O(n8116) );
  INVNHD U7663 ( .I(n12562), .O(n6539) );
  NR2GHD U7664 ( .I1(n11469), .I2(n11470), .O(n11472) );
  ND2KHD U7665 ( .I1(n6729), .I2(n11365), .O(n6540) );
  INVQHD U7666 ( .I(_i_CLEFIA128_keyK _65), .O(n13714) );
  NR2GHD U7667 ( .I1(n11361), .I2(n10054), .O(n7668) );
  ND3EHD U7668 ( .I1(n7025), .I2(n9416), .I3(n12735), .O(n11357) );
  INVCKLHD U7669 ( .I(n6613), .O(n7314) );
  ND2HHD U7670 ( .I1(n6542), .I2(_i_CLEFIA128_keyK _106), .O(n11877) );
  NR2GHD U7671 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(n8798), .O(n6542) );
  INVCKLHD U7672 ( .I(n6666), .O(n7320) );
  OA112HHD U7673 ( .C1(n8792), .C2(n12770), .A1(n9666), .B1(n12768), .O(n12772) );
  NR2IHD U7674 ( .I1(n9332), .I2(n8606), .O(n7105) );
  ND2KHD U7675 ( .I1(n10266), .I2(n9830), .O(n8606) );
  BUFMHD U7676 ( .I(n9918), .O(n9917) );
  ND3EHD U7677 ( .I1(n8495), .I2(n8888), .I3(n10825), .O(n10748) );
  ND2HHD U7678 ( .I1(n12677), .I2(n12688), .O(n10749) );
  ND2HHD U7679 ( .I1(n6544), .I2(n6984), .O(n7406) );
  NR2GHD U7680 ( .I1(n6545), .I2(n12345), .O(n6544) );
  ND2DHD U7681 ( .I1(n12436), .I2(n12361), .O(n6545) );
  ND3EHD U7682 ( .I1(n6546), .I2(n9204), .I3(n9203), .O(n9202) );
  ND3EHD U7683 ( .I1(n9091), .I2(n9201), .I3(n9200), .O(n6546) );
  ND3EHD U7684 ( .I1(n6547), .I2(n10275), .I3(n10038), .O(n9255) );
  NR2GHD U7685 ( .I1(n10274), .I2(n9064), .O(n6547) );
  OA12HHD U7686 ( .B1(n13157), .B2(n13156), .A1(n13634), .O(n13158) );
  NR2IHD U7687 ( .I1(n8153), .I2(n11998), .O(n12118) );
  ND2KHD U7688 ( .I1(n9207), .I2(n9857), .O(n11998) );
  NR2IHD U7689 ( .I1(n9942), .I2(n10807), .O(n11229) );
  NR2IHD U7690 ( .I1(n8902), .I2(n8797), .O(n6779) );
  ND2HHD U7691 ( .I1(n7931), .I2(n7537), .O(n11805) );
  NR2EHD U7692 ( .I1(n13495), .I2(n13238), .O(n7353) );
  ND2HHD U7693 ( .I1(n9831), .I2(n9606), .O(n7129) );
  NR2IHD U7694 ( .I1(n7584), .I2(n7583), .O(n9831) );
  INVKHD U7695 ( .I(n6548), .O(n12172) );
  ND2HHD U7696 ( .I1(n7383), .I2(n11679), .O(n6548) );
  BUFNHD U7697 ( .I(n12264), .O(n8153) );
  NR2IHD U7698 ( .I1(n13809), .I2(n9178), .O(n11730) );
  INVKHD U7699 ( .I(n9887), .O(n8990) );
  NR2IHD U7700 ( .I1(n13184), .I2(n12042), .O(n12398) );
  ND3EHD U7701 ( .I1(n10228), .I2(n10131), .I3(n11996), .O(n7969) );
  OR3HHD U7702 ( .I1(n11434), .I2(n9899), .I3(n9388), .O(n12463) );
  ND2DHD U7703 ( .I1(n11681), .I2(n7538), .O(n8260) );
  ND2HHD U7704 ( .I1(n13175), .I2(n6550), .O(n6549) );
  INVCKGHD U7705 ( .I(n9165), .O(n6550) );
  ND3EHD U7706 ( .I1(n8447), .I2(n10315), .I3(n6851), .O(n10317) );
  ND2KHD U7707 ( .I1(n7051), .I2(_i_CLEFIA128_keyK _120), .O(n11591) );
  ND2KHD U7708 ( .I1(n12905), .I2(n12287), .O(n13150) );
  ND2KHD U7709 ( .I1(n7499), .I2(n11403), .O(n10070) );
  BUFKHD U7710 ( .I(n11677), .O(n6551) );
  INVKHD U7711 ( .I(n6552), .O(n13607) );
  ND3EHD U7712 ( .I1(n12043), .I2(n12398), .I3(n12374), .O(n6552) );
  ND2KHD U7713 ( .I1(n7081), .I2(n6553), .O(n8776) );
  ND2KHD U7714 ( .I1(n11843), .I2(n6840), .O(n9518) );
  ND3EHD U7715 ( .I1(n10592), .I2(n12473), .I3(n11525), .O(n10611) );
  ND2HHD U7716 ( .I1(n8250), .I2(n8420), .O(n10155) );
  NR2GHD U7717 ( .I1(n7702), .I2(n7290), .O(n8420) );
  INVMHD U7718 ( .I(n8187), .O(n6836) );
  ND2HHD U7719 ( .I1(n10739), .I2(n10738), .O(n10755) );
  AN2HHD U7720 ( .I1(n9208), .I2(n12501), .O(n8409) );
  ND2HHD U7721 ( .I1(n7559), .I2(n8290), .O(n7558) );
  NR2GHD U7722 ( .I1(n7804), .I2(n6555), .O(n7802) );
  NR2GHD U7723 ( .I1(n8120), .I2(n13015), .O(n8119) );
  ND2HHD U7724 ( .I1(n6557), .I2(n6556), .O(n8000) );
  INVKHD U7725 ( .I(n6558), .O(n12672) );
  ND2HHD U7726 ( .I1(n8808), .I2(n8807), .O(n6558) );
  NR2CHD U7727 ( .I1(n13619), .I2(n12277), .O(n12278) );
  XNR2KHD U7728 ( .I1(n6821), .I2(n6559), .O(n15067) );
  XOR2HHD U7729 ( .I1(n14214), .I2(n14213), .O(n6559) );
  AN3HHD U7730 ( .I1(n13096), .I2(n13077), .I3(n7842), .O(n9355) );
  ND2KHD U7731 ( .I1(n7292), .I2(n7907), .O(n7842) );
  AN3HHD U7732 ( .I1(n7618), .I2(n7620), .I3(_i_CLEFIA128_state_reg _1), .O(n7878) );
  BUFNHD U7733 ( .I(n12750), .O(n9049) );
  ND2HHD U7734 ( .I1(n13183), .I2(n12401), .O(n12102) );
  BUFEHD U7735 ( .I(n10563), .O(n6560) );
  ND2KHD U7736 ( .I1(n9766), .I2(n9730), .O(n12611) );
  INVLHD U7737 ( .I(n8760), .O(n7291) );
  NR2GHD U7738 ( .I1(n6561), .I2(n9765), .O(n7805) );
  ND3EHD U7739 ( .I1(n9144), .I2(n11546), .I3(n11530), .O(n6561) );
  INVMHD U7740 ( .I(n7046), .O(n8183) );
  ND2KHD U7741 ( .I1(n7280), .I2(n7275), .O(n7274) );
  ND2KHD U7742 ( .I1(n7975), .I2(n6925), .O(n7973) );
  NR2CHD U7743 ( .I1(n13480), .I2(n10002), .O(n9552) );
  OR3HHD U7744 ( .I1(n6650), .I2(n6649), .I3(n9823), .O(n13480) );
  NR2IHD U7745 ( .I1(n10187), .I2(n7699), .O(n7074) );
  INVNHD U7746 ( .I(_i_CLEFIA128_keyL _123), .O(n15074) );
  ND2HHD U7747 ( .I1(n8734), .I2(n8302), .O(n8733) );
  INVDHD U7748 ( .I(n8804), .O(n10824) );
  NR2EHD U7749 ( .I1(n7980), .I2(n7793), .O(n9852) );
  ND3EHD U7750 ( .I1(n6563), .I2(n14055), .I3(n11744), .O(n11651) );
  AN2HHD U7751 ( .I1(n14072), .I2(n13077), .O(n6563) );
  ND3EHD U7752 ( .I1(n6565), .I2(n7681), .I3(n6564), .O(n12557) );
  INVGHD U7753 ( .I(n6861), .O(n6564) );
  INVGHD U7754 ( .I(n8017), .O(n6565) );
  INVCKIHD U7755 ( .I(n6566), .O(n7163) );
  ND3EHD U7756 ( .I1(n12366), .I2(n8887), .I3(n12338), .O(n6566) );
  BUFEHD U7757 ( .I(n7833), .O(n6567) );
  ND2HHD U7758 ( .I1(n10107), .I2(n11929), .O(n8780) );
  NR2IHD U7759 ( .I1(n8126), .I2(n8763), .O(n11929) );
  ND3EHD U7760 ( .I1(n6568), .I2(n7021), .I3(n11322), .O(n10175) );
  ND2KHD U7761 ( .I1(n7656), .I2(n8510), .O(n12576) );
  ND3EHD U7762 ( .I1(n12556), .I2(n6569), .I3(n6922), .O(n7284) );
  NR2EHD U7763 ( .I1(n12757), .I2(n12552), .O(n6569) );
  BUFEHD U7764 ( .I(n14053), .O(n6571) );
  NR2GHD U7765 ( .I1(n13380), .I2(n13379), .O(n13418) );
  ND2HHD U7766 ( .I1(n8515), .I2(n11410), .O(n11352) );
  ND3CHD U7767 ( .I1(n10502), .I2(n9473), .I3(n9470), .O(n9469) );
  INVGHD U7768 ( .I(n6572), .O(n9284) );
  ND2HHD U7769 ( .I1(n7139), .I2(n13035), .O(n6572) );
  ND3CHD U7770 ( .I1(n11526), .I2(n11304), .I3(n11303), .O(n11309) );
  NR2GHD U7771 ( .I1(n12760), .I2(n12759), .O(n12764) );
  AN2HHD U7772 ( .I1(n11296), .I2(n11295), .O(n11298) );
  AN2HHD U7773 ( .I1(n9794), .I2(n14405), .O(n9793) );
  INVGHD U7774 ( .I(n11864), .O(n9586) );
  AN3HHD U7775 ( .I1(n11440), .I2(n11522), .I3(n12486), .O(n7091) );
  INVGHD U7776 ( .I(n10820), .O(n7982) );
  AN2HHD U7777 ( .I1(n13419), .I2(n13420), .O(n6986) );
  NR2EHD U7778 ( .I1(n6876), .I2(n7099), .O(n9843) );
  NR2GHD U7779 ( .I1(n8098), .I2(n8096), .O(n7153) );
  INVGHD U7780 ( .I(n6573), .O(n7366) );
  ND3CHD U7781 ( .I1(n7223), .I2(n7454), .I3(n7340), .O(n6573) );
  OA12HHD U7782 ( .B1(n9895), .B2(n15512), .A1(n8281), .O(n7999) );
  ND2KHD U7783 ( .I1(n8254), .I2(n14055), .O(n13224) );
  ND2KHD U7784 ( .I1(n7362), .I2(n9482), .O(n7150) );
  INVJHD U7785 ( .I(n11614), .O(n11843) );
  NR2IHD U7786 ( .I1(n6823), .I2(n12189), .O(n8079) );
  ND3EHD U7787 ( .I1(n12522), .I2(n10847), .I3(n12619), .O(n6574) );
  ND2KHD U7788 ( .I1(n12619), .I2(n10806), .O(n9942) );
  BUFMHD U7789 ( .I(n8074), .O(n7613) );
  ND3EHD U7790 ( .I1(n12332), .I2(n12331), .I3(n13397), .O(n12333) );
  ND2KHD U7791 ( .I1(n12656), .I2(n11070), .O(n7396) );
  NR2IHD U7792 ( .I1(n10547), .I2(n10548), .O(n7915) );
  ND2HHD U7793 ( .I1(n6580), .I2(n6579), .O(n8045) );
  INVJHD U7794 ( .I(n9494), .O(n6580) );
  NR2IHD U7795 ( .I1(n6581), .I2(n6585), .O(n9558) );
  OA13EHD U7796 ( .B1(n13073), .B2(n13075), .B3(n13074), .A1(n14067), .O(n6581) );
  ND3EHD U7797 ( .I1(n11773), .I2(n12089), .I3(n12298), .O(n11732) );
  ND2HHD U7798 ( .I1(n7809), .I2(n8196), .O(n11773) );
  BUFEHD U7799 ( .I(n13642), .O(n6582) );
  ND3EHD U7800 ( .I1(n6703), .I2(n7162), .I3(n7816), .O(n7813) );
  ND3EHD U7801 ( .I1(n10875), .I2(n11236), .I3(n9145), .O(n10876) );
  ND2KHD U7802 ( .I1(n10011), .I2(n10668), .O(n11236) );
  ND2HHD U7803 ( .I1(n9175), .I2(n9720), .O(n6583) );
  INVGHD U7804 ( .I(n9357), .O(n12207) );
  INVMHD U7805 ( .I(n6584), .O(n8195) );
  NR2IHD U7806 ( .I1(n9333), .I2(n12075), .O(n6584) );
  OR3HHD U7807 ( .I1(n9257), .I2(n12531), .I3(n6813), .O(n12536) );
  INVNHD U7808 ( .I(n9516), .O(n9628) );
  INVJHD U7809 ( .I(n10002), .O(n8149) );
  OA13EHD U7810 ( .B1(n13065), .B2(n13498), .B3(n13064), .A1(n14087), .O(n6585) );
  ND2KHD U7811 ( .I1(n14080), .I2(n8253), .O(n7717) );
  ND2KHD U7812 ( .I1(n6704), .I2(n6735), .O(n7758) );
  NR2IHD U7813 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(n9995), .O(n7762) );
  BUFKHD U7814 ( .I(n8061), .O(n6587) );
  BUFKHD U7815 ( .I(n13098), .O(n6589) );
  ND3EHD U7816 ( .I1(n6590), .I2(n10108), .I3(n10110), .O(n8845) );
  ND2HHD U7817 ( .I1(n11866), .I2(n11874), .O(n6590) );
  ND2KHD U7818 ( .I1(n9038), .I2(n9035), .O(n13767) );
  OA22HHD U7819 ( .A1(n11639), .A2(n11638), .B1(n11658), .B2(n9692), .O(n9038));
  INVCKIHD U7820 ( .I(n8212), .O(n10660) );
  NR2IHD U7821 ( .I1(n9456), .I2(n12133), .O(n11993) );
  ND2KHD U7822 ( .I1(n12120), .I2(n9206), .O(n12133) );
  XOR2HHD U7823 ( .I1(n8787), .I2(n6591), .O(n6662) );
  ND2HHD U7824 ( .I1(n10153), .I2(n13113), .O(n6591) );
  NR2IHD U7825 ( .I1(n9819), .I2(n6592), .O(n9664) );
  ND2HHD U7826 ( .I1(n9112), .I2(n13468), .O(n6592) );
  INVKHD U7827 ( .I(n8213), .O(n8203) );
  ND3EHD U7828 ( .I1(n13596), .I2(n12934), .I3(n13195), .O(n12288) );
  ND2KHD U7829 ( .I1(n8116), .I2(n9050), .O(n12727) );
  INVDHD U7830 ( .I(n9411), .O(n10032) );
  INVDHD U7831 ( .I(DOUT_82), .O(n9947) );
  NR2GHD U7832 ( .I1(n9436), .I2(n12346), .O(n9437) );
  ND3EHD U7833 ( .I1(n8531), .I2(n10423), .I3(n10283), .O(n7589) );
  ND2HHD U7834 ( .I1(n6593), .I2(_i_CLEFIA128_state_reg _1), .O(n7451) );
  ND3EHD U7835 ( .I1(n10407), .I2(n14991), .I3(_i_CLEFIA128_rndcnt_reg _0), .O(n6593) );
  ND3EHD U7836 ( .I1(n6594), .I2(n15176), .I3(_i_CLEFIA128_rndcnt_reg _0), .O(n6614) );
  ND2HHD U7837 ( .I1(n8039), .I2(_i_CLEFIA128_keyK _29), .O(n6594) );
  ND2HHD U7838 ( .I1(n8127), .I2(n11629), .O(n8860) );
  INVKHD U7839 ( .I(n14707), .O(n7433) );
  INVKHD U7840 ( .I(n6595), .O(n9978) );
  ND3EHD U7841 ( .I1(n7802), .I2(n6731), .I3(n7800), .O(n6595) );
  ND2KHD U7842 ( .I1(n12988), .I2(n12361), .O(n9675) );
  ND2KHD U7843 ( .I1(n12226), .I2(n7038), .O(n12361) );
  INVHHD U7844 ( .I(n10836), .O(n6841) );
  AO22HHD U7845 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _116), .B1(n15504), .B2(_i_CLEFIA128_keyK _52), .O(n8286) );
  INVGHD U7846 ( .I(n10549), .O(n10185) );
  INVJHD U7847 ( .I(n12787), .O(n7824) );
  INVHHD U7848 ( .I(n13005), .O(n11936) );
  INVGHD U7849 ( .I(n12793), .O(n8529) );
  INVNHD U7850 ( .I(n10183), .O(n12030) );
  AN3HHD U7851 ( .I1(n11987), .I2(n9322), .I3(n9321), .O(n9320) );
  ND3EHD U7852 ( .I1(n7245), .I2(n6937), .I3(n7594), .O(n7356) );
  NR2IHD U7853 ( .I1(n13489), .I2(n11616), .O(n7245) );
  INVQHD U7854 ( .I(n6599), .O(n7034) );
  INVLHD U7855 ( .I(n8079), .O(n6599) );
  ND3EHD U7856 ( .I1(n6601), .I2(n6600), .I3(n12747), .O(n8865) );
  ND3EHD U7857 ( .I1(n7196), .I2(n8455), .I3(n8682), .O(n6600) );
  ND3EHD U7858 ( .I1(n8457), .I2(n8459), .I3(n12723), .O(n6601) );
  NR2IHD U7859 ( .I1(n10647), .I2(n9331), .O(n10327) );
  INVCKIHD U7860 ( .I(n6602), .O(n6987) );
  ND2HHD U7861 ( .I1(n10855), .I2(n11233), .O(n6602) );
  AN2HHD U7862 ( .I1(n7580), .I2(n9344), .O(n7579) );
  INVJHD U7863 ( .I(n6603), .O(n8904) );
  INVJHD U7864 ( .I(n12750), .O(n6603) );
  AN2HHD U7865 ( .I1(n10791), .I2(n10384), .O(n10023) );
  ND2CHD U7866 ( .I1(n13607), .I2(n8446), .O(n12116) );
  INVJHD U7867 ( .I(n8199), .O(n9330) );
  ND2KHD U7868 ( .I1(n12677), .I2(n10728), .O(n10907) );
  ND3EHD U7869 ( .I1(n9754), .I2(n12979), .I3(n12978), .O(n12980) );
  ND2KHD U7870 ( .I1(n8176), .I2(n7567), .O(n10471) );
  INVJHD U7871 ( .I(n10138), .O(n9412) );
  ND2KHD U7872 ( .I1(n7677), .I2(n7548), .O(n8773) );
  NR2IHD U7873 ( .I1(n7014), .I2(n11505), .O(n7548) );
  ND2KHD U7874 ( .I1(n11070), .I2(n11262), .O(n11212) );
  ND2HHD U7875 ( .I1(n14082), .I2(n11744), .O(n6605) );
  OR3HHD U7876 ( .I1(n13127), .I2(n13126), .I3(n10132), .O(n6606) );
  OAI12CHD U7877 ( .B1(n11960), .B2(n11961), .A1(n13426), .O(n7631) );
  BUFEHD U7878 ( .I(n13460), .O(n6607) );
  ND3EHD U7879 ( .I1(n6608), .I2(_i_CLEFIA128_rndcnt_reg _0), .I3(n15198), .O(n11569) );
  ND2HHD U7880 ( .I1(n6609), .I2(_i_CLEFIA128_keyK _57), .O(n6608) );
  INVCKGHD U7881 ( .I(n8798), .O(n6609) );
  NR2IHD U7882 ( .I1(n11903), .I2(n11911), .O(n11897) );
  NR2GHD U7883 ( .I1(n9361), .I2(n6610), .O(n8640) );
  OR3HHD U7884 ( .I1(n12791), .I2(n12789), .I3(n7476), .O(n6610) );
  ND2KHD U7885 ( .I1(n12656), .I2(n10806), .O(n7177) );
  INVCKLHD U7886 ( .I(n10761), .O(n8859) );
  ND2HHD U7887 ( .I1(n7784), .I2(n9572), .O(n7160) );
  ND3EHD U7888 ( .I1(n12547), .I2(n12545), .I3(n12546), .O(n12548) );
  AOI13BHD U7889 ( .B1(n10524), .B2(n10523), .B3(n12590), .A1(n6611), .O(n7125) );
  INVCKLHD U7890 ( .I(n10426), .O(n10152) );
  ND3EHD U7891 ( .I1(n6612), .I2(n12865), .I3(n12864), .O(n7741) );
  ND2HHD U7892 ( .I1(n7743), .I2(n12855), .O(n6612) );
  INVMHD U7893 ( .I(_i_CLEFIA128_keyL _37), .O(n15047) );
  ND2DHD U7894 ( .I1(n10969), .I2(n8215), .O(n7475) );
  INVGHD U7895 ( .I(n13371), .O(n11955) );
  AN2HHD U7896 ( .I1(n10080), .I2(n13590), .O(n8391) );
  NR2GHD U7897 ( .I1(n12289), .I2(n12288), .O(n12899) );
  NR2IHD U7898 ( .I1(n12377), .I2(n10228), .O(n13593) );
  ND2KHD U7899 ( .I1(n11996), .I2(n10131), .O(n12377) );
  ND3CHD U7900 ( .I1(n8039), .I2(n14817), .I3(_i_CLEFIA128_keyK _107), .O(n11858) );
  NR2IHD U7901 ( .I1(n14152), .I2(n14151), .O(n14153) );
  ND2HHD U7902 ( .I1(n6614), .I2(_i_CLEFIA128_state_reg _1), .O(n6613) );
  INVMHD U7903 ( .I(n6616), .O(n12596) );
  ND2HHD U7904 ( .I1(n9145), .I2(n7365), .O(n6616) );
  BUFEHD U7905 ( .I(n11063), .O(n6617) );
  AN2HHD U7906 ( .I1(n11216), .I2(n11234), .O(n11237) );
  ND2HHD U7907 ( .I1(n11262), .I2(n7359), .O(n10842) );
  NR2IHD U7908 ( .I1(n10842), .I2(n12658), .O(n10846) );
  INVQHD U7909 ( .I(_i_CLEFIA128_keyK _66), .O(n7575) );
  ND3EHD U7910 ( .I1(n7965), .I2(n11828), .I3(n11827), .O(n11837) );
  NR2IHD U7911 ( .I1(n6620), .I2(n6619), .O(n7965) );
  ND2HHD U7912 ( .I1(n6934), .I2(n12198), .O(n6620) );
  NR2IHD U7913 ( .I1(n11242), .I2(n10679), .O(n10680) );
  INVKHD U7914 ( .I(n9078), .O(n10096) );
  BUFEHD U7915 ( .I(n11503), .O(n6621) );
  INVQHD U7916 ( .I(n8798), .O(n6622) );
  INVNHD U7917 ( .I(_i_CLEFIA128_keyK _125), .O(n9498) );
  OAI12CHD U7918 ( .B1(n6623), .B2(n9419), .A1(n8498), .O(n8035) );
  NR2GHD U7919 ( .I1(n7224), .I2(n14707), .O(n6623) );
  INVDHD U7920 ( .I(n6728), .O(n6727) );
  ND3EHD U7921 ( .I1(n11377), .I2(n11371), .I3(n11105), .O(n11106) );
  NR2EHD U7922 ( .I1(n12941), .I2(n8890), .O(n9981) );
  ND3EHD U7923 ( .I1(n6624), .I2(n11561), .I3(n9497), .O(n11564) );
  AN2HHD U7924 ( .I1(n11562), .I2(n14405), .O(n6624) );
  ND2HHD U7925 ( .I1(n6820), .I2(n12731), .O(n11102) );
  ND2KHD U7926 ( .I1(n9209), .I2(n7015), .O(n10619) );
  INVKHD U7927 ( .I(n8218), .O(n6882) );
  ND2HHD U7928 ( .I1(n6625), .I2(n6626), .O(n11582) );
  OA112HHD U7929 ( .C1(n11581), .C2(n11580), .A1(n11579), .B1(_i_CLEFIA128_state_reg _1), .O(n6625) );
  ND3EHD U7930 ( .I1(n11578), .I2(n11577), .I3(n11576), .O(n6626) );
  XOR2HHD U7931 ( .I1(n8948), .I2(n6627), .O(n7225) );
  ND3EHD U7932 ( .I1(n7226), .I2(n7096), .I3(n8687), .O(n6627) );
  INVKHD U7933 ( .I(n12878), .O(n7030) );
  INVGHD U7934 ( .I(n13251), .O(n6628) );
  ND2HHD U7935 ( .I1(n7044), .I2(n6628), .O(n8358) );
  ND2KHD U7936 ( .I1(_i_CLEFIA128_keyK _88), .I2(n8797), .O(n8497) );
  NR2IHD U7937 ( .I1(n6833), .I2(n11021), .O(n11334) );
  ND2KHD U7938 ( .I1(n10259), .I2(n9840), .O(n11021) );
  ND2HHD U7939 ( .I1(n6631), .I2(n6630), .O(n10590) );
  INVCKGHD U7940 ( .I(n11300), .O(n6630) );
  XNR2HHD U7941 ( .I1(n10582), .I2(n10581), .O(n11300) );
  ND3EHD U7942 ( .I1(n11402), .I2(n10073), .I3(n7307), .O(n7098) );
  ND2HHD U7943 ( .I1(n9964), .I2(n11176), .O(n9615) );
  INVJHD U7944 ( .I(n12475), .O(n6855) );
  BUFEHD U7945 ( .I(n13216), .O(n6632) );
  ND2HHD U7946 ( .I1(n7667), .I2(n11479), .O(n7666) );
  ND2HHD U7947 ( .I1(n13801), .I2(n13800), .O(n6096) );
  NR2EHD U7948 ( .I1(n10627), .I2(n10694), .O(n10629) );
  ND2HHD U7949 ( .I1(n13036), .I2(n9574), .O(n12340) );
  INVGHD U7950 ( .I(n6633), .O(n12253) );
  ND2HHD U7951 ( .I1(n12252), .I2(n13460), .O(n6633) );
  ND3EHD U7952 ( .I1(n12743), .I2(n6820), .I3(n11349), .O(n10515) );
  ND3EHD U7953 ( .I1(n7060), .I2(n7062), .I3(n6634), .O(n7387) );
  XOR2HHD U7954 ( .I1(n14168), .I2(n8031), .O(n13961) );
  XOR2HHD U7955 ( .I1(n13767), .I2(n7943), .O(n10218) );
  ND2KHD U7956 ( .I1(n7838), .I2(n9803), .O(n7943) );
  OR3HHD U7957 ( .I1(n8015), .I2(n11321), .I3(n12738), .O(n12592) );
  XNR2KHD U7958 ( .I1(n9930), .I2(n13557), .O(n14913) );
  INVKHD U7959 ( .I(n7664), .O(n7662) );
  ND3EHD U7960 ( .I1(n9391), .I2(n15306), .I3(_i_CLEFIA128_rndcnt_reg _0), .O(n8999) );
  NR2GHD U7961 ( .I1(n12348), .I2(n9404), .O(n9301) );
  BUFMHD U7962 ( .I(n10481), .O(n9099) );
  ND2KHD U7963 ( .I1(n8895), .I2(n7917), .O(n8796) );
  NR2IHD U7964 ( .I1(n10213), .I2(n10055), .O(n8895) );
  INVMHD U7965 ( .I(n6931), .O(n11679) );
  BUFEHD U7966 ( .I(n9873), .O(n6635) );
  INVKHD U7967 ( .I(n9505), .O(n13232) );
  INVGHD U7968 ( .I(n12208), .O(n8148) );
  ND3EHD U7969 ( .I1(n8951), .I2(n8950), .I3(n8949), .O(n6636) );
  INVKHD U7970 ( .I(n12537), .O(n10877) );
  ND3EHD U7971 ( .I1(n6638), .I2(n8342), .I3(n6637), .O(n6169) );
  ND2HHD U7972 ( .I1(n6887), .I2(n15500), .O(n6637) );
  NR2EHD U7973 ( .I1(n11807), .I2(n7861), .O(n11808) );
  BUFNHD U7974 ( .I(n9731), .O(n7161) );
  BUFKHD U7975 ( .I(n14059), .O(n6639) );
  NR2IHD U7976 ( .I1(n10658), .I2(n10657), .O(n10664) );
  ND2HHD U7977 ( .I1(n14080), .I2(n7118), .O(n6640) );
  ND2KHD U7978 ( .I1(n9547), .I2(n9041), .O(n8755) );
  AN2HHD U7979 ( .I1(n12917), .I2(n8657), .O(n8656) );
  AN3HHD U7980 ( .I1(n8638), .I2(n8634), .I3(n8636), .O(n8984) );
  ND2DHD U7981 ( .I1(n10315), .I2(n7389), .O(n10316) );
  AO22HHD U7982 ( .A1(n7045), .A2(n13256), .B1(n15504), .B2(n13255), .O(n10290) );
  XNR2KHD U7983 ( .I1(_i_CLEFIA128_CON_T_x _3), .I2(DOUT_42), .O(n8975) );
  AN2HHD U7984 ( .I1(_i_CLEFIA128_keyK _48), .I2(_i_CLEFIA128_keyL _48), .O(n8379) );
  NR2EHD U7985 ( .I1(n6642), .I2(n13136), .O(n13138) );
  ND3EHD U7986 ( .I1(n13131), .I2(n13130), .I3(n7165), .O(n6642) );
  AN2HHD U7987 ( .I1(n11737), .I2(n11736), .O(n8294) );
  ND2HHD U7988 ( .I1(n9898), .I2(n11018), .O(n11410) );
  ND2HHD U7989 ( .I1(n10215), .I2(n9539), .O(n9971) );
  NR2EHD U7990 ( .I1(n12803), .I2(n12802), .O(n12804) );
  ND2KHD U7991 ( .I1(n7035), .I2(n7254), .O(n12087) );
  NR2GHD U7992 ( .I1(n11352), .I2(n11351), .O(n11353) );
  AN3HHD U7993 ( .I1(n8420), .I2(n8221), .I3(n8253), .O(n13057) );
  XOR2HHD U7994 ( .I1(n14328), .I2(n14329), .O(n10161) );
  ND2HHD U7995 ( .I1(n9046), .I2(n11856), .O(n14328) );
  XNR2KHD U7996 ( .I1(n13767), .I2(n7943), .O(n10149) );
  ND3EHD U7997 ( .I1(n6705), .I2(n13072), .I3(n12197), .O(n7910) );
  INVNHD U7998 ( .I(n7865), .O(n10802) );
  BUFEHD U7999 ( .I(n12669), .O(n6643) );
  ND2HHD U8000 ( .I1(n11787), .I2(n7537), .O(n6644) );
  NR2EHD U8001 ( .I1(n11651), .I2(n8596), .O(n11656) );
  ND2HHD U8002 ( .I1(n13851), .I2(n13850), .O(n7439) );
  NR2IHD U8003 ( .I1(n8058), .I2(n7909), .O(n13851) );
  ND3EHD U8004 ( .I1(n9573), .I2(n7323), .I3(n7834), .O(n10050) );
  ND2HHD U8005 ( .I1(n8743), .I2(_i_CLEFIA128_rndcnt_reg _0), .O(n8742) );
  AN3HHD U8006 ( .I1(n6646), .I2(n7645), .I3(_i_CLEFIA128_state_reg _1), .O(n6778) );
  ND3EHD U8007 ( .I1(n9883), .I2(n15058), .I3(_i_CLEFIA128_rndcnt_reg _0), .O(n6646) );
  OR2HHD U8008 ( .I1(n11087), .I2(n7179), .O(n11088) );
  NR2IHD U8009 ( .I1(n7760), .I2(n7762), .O(n6735) );
  ND3EHD U8010 ( .I1(n12120), .I2(n9206), .I3(n9456), .O(n9635) );
  ND2KHD U8011 ( .I1(n9192), .I2(n10549), .O(n6902) );
  NR2IHD U8012 ( .I1(n11984), .I2(n14707), .O(n9324) );
  INVMHD U8013 ( .I(n7865), .O(n6842) );
  INVQHD U8014 ( .I(_i_CLEFIA128_keyK _121), .O(n8081) );
  ND2HHD U8015 ( .I1(n8797), .I2(_i_CLEFIA128_keyK _1), .O(n10461) );
  NR2IHD U8016 ( .I1(n8207), .I2(n8526), .O(n10424) );
  ND2KHD U8017 ( .I1(n10442), .I2(n10767), .O(n8526) );
  NR2GHD U8018 ( .I1(n7234), .I2(n7233), .O(n8951) );
  ND2KHD U8019 ( .I1(n12651), .I2(n7779), .O(n7346) );
  INVNHD U8020 ( .I(n10091), .O(n10767) );
  ND2KHD U8021 ( .I1(n8927), .I2(n10199), .O(n10202) );
  ND2KHD U8022 ( .I1(n6777), .I2(n6851), .O(n10415) );
  INVQHD U8023 ( .I(n9749), .O(n10746) );
  ND2KHD U8024 ( .I1(n8895), .I2(n7917), .O(n6874) );
  NR2IHD U8025 ( .I1(n11612), .I2(n7500), .O(n8226) );
  ND2KHD U8026 ( .I1(n7977), .I2(n11628), .O(n7500) );
  NR2EHD U8027 ( .I1(n10787), .I2(n10788), .O(n10790) );
  NR2GHD U8028 ( .I1(n8623), .I2(n12300), .O(n8622) );
  NR2IHD U8029 ( .I1(n8117), .I2(n9451), .O(n7489) );
  ND2HHD U8030 ( .I1(n11440), .I2(n12450), .O(n11132) );
  ND2KHD U8031 ( .I1(n9194), .I2(n12498), .O(n12450) );
  ND3EHD U8032 ( .I1(n13099), .I2(n8190), .I3(n12208), .O(n6649) );
  ND2HHD U8033 ( .I1(n13076), .I2(n14071), .O(n6650) );
  NR2IHD U8034 ( .I1(n8883), .I2(n9000), .O(n9804) );
  AN3HHD U8035 ( .I1(n9176), .I2(n8333), .I3(n13814), .O(n8361) );
  NR2GHD U8036 ( .I1(n13514), .I2(n7862), .O(n9176) );
  INVCKGHD U8037 ( .I(n6652), .O(n6651) );
  ND2HHD U8038 ( .I1(n9398), .I2(n13004), .O(n6652) );
  INVCKGHD U8039 ( .I(n6654), .O(n6653) );
  ND2HHD U8040 ( .I1(n9873), .I2(n13036), .O(n6654) );
  NR2IHD U8041 ( .I1(n11671), .I2(n14707), .O(n7578) );
  AN2HHD U8042 ( .I1(n11253), .I2(n9145), .O(n8407) );
  INVNHD U8043 ( .I(n7337), .O(n8315) );
  INVCKIHD U8044 ( .I(n10563), .O(n7619) );
  NR2IHD U8045 ( .I1(n6712), .I2(n8414), .O(n9369) );
  AN2HHD U8046 ( .I1(n8476), .I2(n11091), .O(n8510) );
  INVMHD U8047 ( .I(n8871), .O(n12125) );
  ND2HHD U8048 ( .I1(n7124), .I2(n7123), .O(n12434) );
  NR2EHD U8049 ( .I1(n13631), .I2(n8600), .O(n7950) );
  OR3HHD U8050 ( .I1(n11136), .I2(n11135), .I3(n11134), .O(n11138) );
  AN2HHD U8051 ( .I1(n13661), .I2(n7449), .O(n6962) );
  INVNHD U8052 ( .I(n7833), .O(n9087) );
  ND2KHD U8053 ( .I1(n10619), .I2(n7081), .O(n7833) );
  ND2KHD U8054 ( .I1(n8797), .I2(_i_CLEFIA128_keyK _124), .O(n11586) );
  ND2DHD U8055 ( .I1(n7034), .I2(n13100), .O(n11739) );
  ND2HHD U8056 ( .I1(n8798), .I2(_i_CLEFIA128_keyL _125), .O(n11562) );
  OR2KHD U8057 ( .I1(n11804), .I2(n11710), .O(n8582) );
  INVHHD U8058 ( .I(_i_CLEFIA128_keyL _77), .O(n7349) );
  ND2DHD U8059 ( .I1(n7537), .I2(n13512), .O(n11717) );
  ND2HHD U8060 ( .I1(n7770), .I2(n7771), .O(n7233) );
  ND3EHD U8061 ( .I1(n10526), .I2(n12729), .I3(n6820), .O(n10527) );
  ND3EHD U8062 ( .I1(n6656), .I2(n6655), .I3(n13673), .O(n8835) );
  NR2GHD U8063 ( .I1(n8844), .I2(n11817), .O(n13673) );
  NR3BHD U8064 ( .I1(n8839), .I2(n8842), .I3(n11815), .O(n6655) );
  INVCKGHD U8065 ( .I(n8836), .O(n6656) );
  ND2DHD U8066 ( .I1(n10798), .I2(n7580), .O(n10781) );
  ND2KHD U8067 ( .I1(n10794), .I2(n7507), .O(n7580) );
  ND3EHD U8068 ( .I1(n6657), .I2(n12384), .I3(n6897), .O(n9614) );
  INVCKIHD U8069 ( .I(n6658), .O(n6657) );
  ND2HHD U8070 ( .I1(n9832), .I2(n12935), .O(n6658) );
  ND3EHD U8071 ( .I1(n13812), .I2(n11773), .I3(n13837), .O(n9833) );
  INVMHD U8072 ( .I(n11996), .O(n12913) );
  INVGHD U8073 ( .I(n6659), .O(n12389) );
  ND3EHD U8074 ( .I1(n13199), .I2(n12402), .I3(n8657), .O(n6659) );
  INVGHD U8075 ( .I(n13624), .O(n9039) );
  ND3EHD U8076 ( .I1(n12131), .I2(n12132), .I3(n13211), .O(n13624) );
  NR2GHD U8077 ( .I1(n12161), .I2(n12160), .O(n12166) );
  ND3EHD U8078 ( .I1(n9418), .I2(n14556), .I3(_i_CLEFIA128_rndcnt_reg _0), .O(n7435) );
  ND2KHD U8079 ( .I1(n6660), .I2(n8443), .O(n13615) );
  INVCKIHD U8080 ( .I(n6661), .O(n6660) );
  ND2HHD U8081 ( .I1(n13128), .I2(n13572), .O(n6661) );
  NR2IHD U8082 ( .I1(n10322), .I2(n14707), .O(n9948) );
  ND2KHD U8083 ( .I1(n6615), .I2(n7318), .O(n11062) );
  OA12EHD U8084 ( .B1(n15499), .B2(n15043), .A1(n14669), .O(n8301) );
  BUFCKKHD U8085 ( .I(n13972), .O(n7789) );
  INVNHD U8086 ( .I(n8212), .O(n7863) );
  NR2IHD U8087 ( .I1(n9596), .I2(n13615), .O(n9677) );
  ND3EHD U8088 ( .I1(n11232), .I2(n11231), .I3(n7508), .O(n11247) );
  ND3HHD U8089 ( .I1(n11227), .I2(n11226), .I3(n11225), .O(n11228) );
  INVMHD U8090 ( .I(n12913), .O(n9187) );
  XOR2HHD U8091 ( .I1(n6663), .I2(n6662), .O(n14705) );
  XOR2HHD U8092 ( .I1(n6577), .I2(n14352), .O(n6663) );
  INVLHD U8093 ( .I(n8154), .O(n9206) );
  ND3CHD U8094 ( .I1(n8437), .I2(n11965), .I3(n6796), .O(n9983) );
  NR2EHD U8095 ( .I1(n12597), .I2(n8334), .O(n12602) );
  NR2IHD U8096 ( .I1(n8043), .I2(n8042), .O(n8041) );
  ND2KHD U8097 ( .I1(n11226), .I2(n10806), .O(n11205) );
  ND2KHD U8098 ( .I1(n6842), .I2(n9766), .O(n11226) );
  ND3EHD U8099 ( .I1(n10770), .I2(n9145), .I3(n7580), .O(n10771) );
  ND2HHD U8100 ( .I1(n6665), .I2(n9647), .O(n9075) );
  OA13EHD U8101 ( .B1(n10611), .B2(n11153), .B3(n11310), .A1(n11318), .O(n6665) );
  ND3EHD U8102 ( .I1(n7157), .I2(n6994), .I3(n11219), .O(n10808) );
  ND3EHD U8103 ( .I1(n9584), .I2(n12546), .I3(n9583), .O(n10049) );
  ND2HHD U8104 ( .I1(n10783), .I2(n11063), .O(n6666) );
  INVMHD U8105 ( .I(n8629), .O(n11896) );
  INVGHD U8106 ( .I(n13636), .O(n7951) );
  ND3EHD U8107 ( .I1(n12106), .I2(n8324), .I3(n12105), .O(n13636) );
  ND2HHD U8108 ( .I1(n7940), .I2(n8299), .O(n7939) );
  INVLHD U8109 ( .I(n6818), .O(n6820) );
  NR2GHD U8110 ( .I1(n6668), .I2(n10234), .O(n9397) );
  ND3EHD U8111 ( .I1(n11077), .I2(n12604), .I3(n11217), .O(n6668) );
  ND2HHD U8112 ( .I1(n6778), .I2(n6669), .O(n8747) );
  ND2HHD U8113 ( .I1(n6799), .I2(n11968), .O(n6669) );
  INVJHD U8114 ( .I(n9765), .O(n8782) );
  BUFEHD U8115 ( .I(n12867), .O(n6670) );
  ND3EHD U8116 ( .I1(n12910), .I2(n6918), .I3(n11994), .O(n12026) );
  INVCKGHD U8117 ( .I(n11644), .O(n14057) );
  ND2KHD U8118 ( .I1(n12423), .I2(n9449), .O(n13420) );
  INVGHD U8119 ( .I(n8831), .O(n12158) );
  ND3EHD U8120 ( .I1(n13433), .I2(n9846), .I3(n9342), .O(n13434) );
  NR2GHD U8121 ( .I1(n11754), .I2(n8829), .O(n8072) );
  ND2KHD U8122 ( .I1(n7254), .I2(n8178), .O(n8758) );
  ND2HHD U8123 ( .I1(n12217), .I2(n8234), .O(n9707) );
  AN3HHD U8124 ( .I1(n9679), .I2(n9693), .I3(n12999), .O(n8234) );
  NR2IHD U8125 ( .I1(n10167), .I2(n6759), .O(n9934) );
  AN2HHD U8126 ( .I1(n15263), .I2(_i_CLEFIA128_rndcnt_reg _0), .O(n8370) );
  ND2HHD U8127 ( .I1(n13122), .I2(n8729), .O(n12103) );
  INVGHD U8128 ( .I(n6733), .O(n6732) );
  ND2HHD U8129 ( .I1(n8202), .I2(n9145), .O(n11076) );
  ND2KHD U8130 ( .I1(n6842), .I2(n7864), .O(n8202) );
  BUFEHD U8131 ( .I(n12522), .O(n6671) );
  NR2GHD U8132 ( .I1(n13618), .I2(n13150), .O(n12043) );
  ND3EHD U8133 ( .I1(n12611), .I2(n7185), .I3(n9191), .O(n6673) );
  ND2KHD U8134 ( .I1(n7217), .I2(n9766), .O(n7185) );
  ND2HHD U8135 ( .I1(n9435), .I2(n7933), .O(n9210) );
  ND3EHD U8136 ( .I1(n6674), .I2(n9054), .I3(n9425), .O(n9424) );
  NR2EHD U8137 ( .I1(n9004), .I2(n9005), .O(n6674) );
  INVKHD U8138 ( .I(n12655), .O(n10801) );
  ND2KHD U8139 ( .I1(n10179), .I2(n10178), .O(n12655) );
  ND2HHD U8140 ( .I1(n8525), .I2(n7289), .O(n8524) );
  BUFEHD U8141 ( .I(n12484), .O(n6675) );
  NR2IHD U8142 ( .I1(n12120), .I2(n11998), .O(n11999) );
  NR2EHD U8143 ( .I1(n11238), .I2(n11239), .O(n11244) );
  ND2KHD U8144 ( .I1(n9423), .I2(n7359), .O(n11066) );
  INVLHD U8145 ( .I(n7933), .O(n8006) );
  INVMHD U8146 ( .I(n11905), .O(n10209) );
  INVMHD U8147 ( .I(n10023), .O(n12640) );
  INVJHD U8148 ( .I(n6678), .O(n6869) );
  ND3EHD U8149 ( .I1(n8742), .I2(_i_CLEFIA128_state_reg _1), .I3(n8745), .O(n6678) );
  INVGHD U8150 ( .I(n12435), .O(n12438) );
  ND2DHD U8151 ( .I1(n12637), .I2(n7779), .O(n10835) );
  AN2HHD U8152 ( .I1(n7580), .I2(n12609), .O(n12612) );
  AN2HHD U8153 ( .I1(n8738), .I2(_i_CLEFIA128_rndcnt_reg _0), .O(n7401) );
  ND2HHD U8154 ( .I1(n10388), .I2(n6679), .O(n7602) );
  OAI22CHD U8155 ( .A1(n10382), .A2(n10381), .B1(n10380), .B2(n10379), .O(n6679) );
  INVGHD U8156 ( .I(n11453), .O(n11454) );
  ND3CHD U8157 ( .I1(n11063), .I2(n9145), .I3(n10850), .O(n9027) );
  ND2KHD U8158 ( .I1(n9659), .I2(n10178), .O(n11063) );
  ND2HHD U8159 ( .I1(n7987), .I2(n11663), .O(n6681) );
  INVNHD U8160 ( .I(n8776), .O(n12484) );
  NR2IHD U8161 ( .I1(n12716), .I2(n12667), .O(n9560) );
  ND2KHD U8162 ( .I1(n6931), .I2(n11707), .O(n11775) );
  ND2HHD U8163 ( .I1(n8797), .I2(_i_CLEFIA128_keyK _28), .O(n10310) );
  INVGHD U8164 ( .I(n8511), .O(n12666) );
  ND2HHD U8165 ( .I1(n9785), .I2(n9784), .O(n14015) );
  ND2KHD U8166 ( .I1(n9033), .I2(n11345), .O(n9784) );
  INVGHD U8167 ( .I(n6683), .O(n8820) );
  ND2HHD U8168 ( .I1(n12304), .I2(n13526), .O(n6683) );
  ND2HHD U8169 ( .I1(n7249), .I2(n7248), .O(n10253) );
  INVNHD U8170 ( .I(_i_CLEFIA128_keyL _48), .O(n7251) );
  ND2HHD U8171 ( .I1(n12087), .I2(n9741), .O(n11731) );
  ND2KHD U8172 ( .I1(n10178), .I2(n7507), .O(n7359) );
  ND2KHD U8173 ( .I1(n8577), .I2(n10253), .O(n7416) );
  ND2KHD U8174 ( .I1(n10178), .I2(n6883), .O(n12622) );
  ND3EHD U8175 ( .I1(n11237), .I2(n11235), .I3(n11236), .O(n11238) );
  NR2IHD U8176 ( .I1(n9724), .I2(n11363), .O(n9785) );
  NR2GHD U8177 ( .I1(n13547), .I2(n8085), .O(n7431) );
  BUFEHD U8178 ( .I(n13646), .O(n6685) );
  ND2HHD U8179 ( .I1(n9295), .I2(n7900), .O(n9294) );
  XNR2KHD U8180 ( .I1(_i_CLEFIA128_CON_T_x _9), .I2(DOUT_120), .O(n6925) );
  ND2KHD U8181 ( .I1(n7291), .I2(n7292), .O(n14071) );
  NR2EHD U8182 ( .I1(_i_CLEFIA128_keyK _68), .I2(n14931), .O(n8882) );
  NR2EHD U8183 ( .I1(n7997), .I2(n7996), .O(n7995) );
  INVGHD U8184 ( .I(n11401), .O(n9011) );
  BUFNHD U8185 ( .I(n9802), .O(n7014) );
  ND2HHD U8186 ( .I1(n11119), .I2(n6687), .O(n7685) );
  ND3EHD U8187 ( .I1(n11411), .I2(n7309), .I3(n11511), .O(n6688) );
  INVNHD U8188 ( .I(n7547), .O(n11505) );
  AOI22HHD U8189 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _76), .B1(n15504), .B2(_i_CLEFIA128_keyK _12), .O(n12887) );
  NR2IHD U8190 ( .I1(n11585), .I2(n14707), .O(n9891) );
  NR2IHD U8191 ( .I1(n7674), .I2(n7361), .O(n10512) );
  INVJHD U8192 ( .I(n6689), .O(n8102) );
  ND2KHD U8193 ( .I1(n8797), .I2(_i_CLEFIA128_keyK _0), .O(n6689) );
  NR2GHD U8194 ( .I1(n11092), .I2(n7029), .O(n8476) );
  ND2KHD U8195 ( .I1(n12553), .I2(n8607), .O(n7709) );
  INVQHD U8196 ( .I(_i_CLEFIA128_rndcnt_reg _0), .O(n14405) );
  NR2GHD U8197 ( .I1(n7654), .I2(n7566), .O(n7653) );
  INVGHD U8198 ( .I(n6690), .O(n8280) );
  ND3EHD U8199 ( .I1(n8236), .I2(n10759), .I3(n12866), .O(n6690) );
  ND2KHD U8200 ( .I1(n9162), .I2(n9022), .O(n14140) );
  NR2IHD U8201 ( .I1(n9163), .I2(n9164), .O(n9162) );
  OA12HHD U8202 ( .B1(n6692), .B2(n13094), .A1(n14049), .O(n7300) );
  ND2HHD U8203 ( .I1(n6771), .I2(n14075), .O(n6692) );
  AN2KHD U8204 ( .I1(n7703), .I2(n7336), .O(n7334) );
  ND2KHD U8205 ( .I1(n9194), .I2(n11176), .O(n11297) );
  NR2IHD U8206 ( .I1(n10619), .I2(n10695), .O(n10721) );
  ND2KHD U8207 ( .I1(n9129), .I2(n10587), .O(n10695) );
  ND2KHD U8208 ( .I1(n7051), .I2(_i_CLEFIA128_keyK _98), .O(n11983) );
  ND3EHD U8209 ( .I1(n11641), .I2(n6940), .I3(n6589), .O(n11642) );
  INVCKIHD U8210 ( .I(n10888), .O(n10732) );
  OR3HHD U8211 ( .I1(n13654), .I2(n12168), .I3(n7993), .O(n7992) );
  AN2HHD U8212 ( .I1(n12737), .I2(n11507), .O(n6863) );
  ND2HHD U8213 ( .I1(n8039), .I2(_i_CLEFIA128_keyK _13), .O(n10412) );
  ND2HHD U8214 ( .I1(n6693), .I2(n9312), .O(n13247) );
  NR2GHD U8215 ( .I1(n9314), .I2(n9315), .O(n6693) );
  ND2HHD U8216 ( .I1(n14140), .I2(n14139), .O(n9160) );
  INVMHD U8217 ( .I(n6860), .O(n12423) );
  ND2KHD U8218 ( .I1(n8872), .I2(n11988), .O(n8692) );
  INVLHD U8219 ( .I(n8845), .O(n10107) );
  NR2GHD U8220 ( .I1(n10259), .I2(n6833), .O(n7718) );
  XOR2HHD U8221 ( .I1(_i_CLEFIA128_CON_T_xi _9), .I2(DOUT_34), .O(n10469) );
  ND2HHD U8222 ( .I1(n6696), .I2(n6695), .O(n7628) );
  INVJHD U8223 ( .I(n12357), .O(n6696) );
  ND3CHD U8224 ( .I1(n11981), .I2(n6834), .I3(n6796), .O(n8156) );
  ND2KHD U8225 ( .I1(n10442), .I2(n10091), .O(n9444) );
  ND2HHD U8226 ( .I1(n9462), .I2(n9667), .O(n6697) );
  ND2HHD U8227 ( .I1(n14052), .I2(n7842), .O(n13060) );
  INVGHD U8228 ( .I(n6698), .O(n10730) );
  ND2HHD U8229 ( .I1(n7247), .I2(n10818), .O(n6698) );
  AN2HHD U8230 ( .I1(n11802), .I2(n7687), .O(n6912) );
  ND3EHD U8231 ( .I1(n13182), .I2(n13573), .I3(n13130), .O(n12098) );
  NR2GHD U8232 ( .I1(n9454), .I2(n10951), .O(n10954) );
  ND3EHD U8233 ( .I1(n8664), .I2(_i_CLEFIA128_keyL _113), .I3(n8589), .O(n8663) );
  ND3EHD U8234 ( .I1(n10885), .I2(n8398), .I3(n8921), .O(n9640) );
  AN2HHD U8235 ( .I1(n6970), .I2(n8495), .O(n10885) );
  OR3HHD U8236 ( .I1(n7423), .I2(n6701), .I3(n14068), .O(n8056) );
  OR3HHD U8237 ( .I1(n12186), .I2(n12195), .I3(n12187), .O(n6701) );
  ND2HHD U8238 ( .I1(n8613), .I2(n13492), .O(n11638) );
  NR2GHD U8239 ( .I1(n11613), .I2(n7356), .O(n8613) );
  ND2HHD U8240 ( .I1(n6702), .I2(_i_CLEFIA128_state_reg _1), .O(n8616) );
  ND3EHD U8241 ( .I1(n10412), .I2(n15242), .I3(_i_CLEFIA128_rndcnt_reg _0), .O(n6702) );
  ND3EHD U8242 ( .I1(n7822), .I2(n7820), .I3(n12718), .O(n6703) );
  AN3HHD U8243 ( .I1(n9996), .I2(n11569), .I3(_i_CLEFIA128_state_reg _1), .O(n6704) );
  OR3HHD U8244 ( .I1(n11748), .I2(n10156), .I3(n10155), .O(n8828) );
  ND3EHD U8245 ( .I1(n8548), .I2(n10897), .I3(n12805), .O(n7525) );
  NR2IHD U8246 ( .I1(n10734), .I2(n10733), .O(n12805) );
  OR3HHD U8247 ( .I1(n7717), .I2(n8150), .I3(n7716), .O(n10002) );
  ND2HHD U8248 ( .I1(n7452), .I2(n9448), .O(n7242) );
  NR2IHD U8249 ( .I1(n8560), .I2(n8559), .O(n7452) );
  XNR2KHD U8250 ( .I1(n14171), .I2(n7381), .O(n6787) );
  XNR2KHD U8251 ( .I1(n10019), .I2(n10020), .O(n14633) );
  ND2KHD U8252 ( .I1(n9615), .I2(n9135), .O(n9446) );
  OR2KHD U8253 ( .I1(n9989), .I2(n11863), .O(n9268) );
  OA13EHD U8254 ( .B1(n12444), .B2(n7484), .B3(n8625), .A1(n13426), .O(n9861));
  ND3EHD U8255 ( .I1(n12438), .I2(n8119), .I3(n12437), .O(n7484) );
  ND2HHD U8256 ( .I1(n8434), .I2(n6708), .O(n8551) );
  INVCKGHD U8257 ( .I(n8798), .O(n6709) );
  ND2HHD U8258 ( .I1(n7487), .I2(n9693), .O(n8120) );
  ND3CHD U8259 ( .I1(n6710), .I2(n8588), .I3(n14405), .O(n7781) );
  ND3EHD U8260 ( .I1(n15189), .I2(n8797), .I3(_i_CLEFIA128_keyK _72), .O(n6710) );
  ND3EHD U8261 ( .I1(n7888), .I2(n7887), .I3(n6916), .O(n7882) );
  AN2HHD U8262 ( .I1(n12668), .I2(n7340), .O(n6916) );
  ND3EHD U8263 ( .I1(n11484), .I2(n8484), .I3(n9619), .O(n11107) );
  NR2IHD U8264 ( .I1(n7720), .I2(n8134), .O(n9431) );
  ND2KHD U8265 ( .I1(n7783), .I2(n9431), .O(n8778) );
  NR2IHD U8266 ( .I1(n10209), .I2(n12216), .O(n8851) );
  ND3EHD U8267 ( .I1(n14054), .I2(n6571), .I3(n14052), .O(n14064) );
  ND2HHD U8268 ( .I1(n10550), .I2(n7389), .O(n9192) );
  ND2HHD U8269 ( .I1(n10005), .I2(n13122), .O(n12255) );
  ND3EHD U8270 ( .I1(n7139), .I2(n13425), .I3(n8392), .O(n12218) );
  ND3CHD U8271 ( .I1(n8039), .I2(n8982), .I3(_i_CLEFIA128_keyK _101), .O(n11971) );
  XOR2HHD U8272 ( .I1(_i_CLEFIA128_keyL _122), .I2(n11573), .O(n11575) );
  INVCKGHD U8273 ( .I(n13438), .O(n13456) );
  XOR2HHD U8274 ( .I1(n13556), .I2(n14993), .O(n14364) );
  NR2GHD U8275 ( .I1(n12185), .I2(n8860), .O(n11633) );
  INVKHD U8276 ( .I(n10446), .O(n8134) );
  NR2GHD U8277 ( .I1(n13230), .I2(n8829), .O(n13240) );
  XNR2KHD U8278 ( .I1(_i_CLEFIA128_keyL _93), .I2(n8174), .O(n10315) );
  OA13EHD U8279 ( .B1(n13485), .B2(n13484), .B3(n13486), .A1(n14087), .O(n6712) );
  NR2GHD U8280 ( .I1(n10769), .I2(n10766), .O(n8494) );
  OA12HHD U8281 ( .B1(n10008), .B2(n11129), .A1(n14808), .O(n7902) );
  ND2KHD U8282 ( .I1(n11402), .I2(n10534), .O(n9086) );
  ND3EHD U8283 ( .I1(n8944), .I2(n15352), .I3(_i_CLEFIA128_rndcnt_reg _0), .O(n7228) );
  ND2KHD U8284 ( .I1(_i_CLEFIA128_keyK _9), .I2(n8797), .O(n8944) );
  ND3EHD U8285 ( .I1(n9053), .I2(n10625), .I3(n12450), .O(n10626) );
  XOR2HHD U8286 ( .I1(n9962), .I2(n6713), .O(n9151) );
  XOR2HHD U8287 ( .I1(n14804), .I2(n13952), .O(n6713) );
  ND2KHD U8288 ( .I1(n9898), .I2(n9694), .O(n12558) );
  ND3EHD U8289 ( .I1(n10188), .I2(n7389), .I3(n11575), .O(n8024) );
  XNR2KHD U8290 ( .I1(DOUT_58), .I2(_i_CLEFIA128_CON_T_xi _9), .O(n9411) );
  ND2HHD U8291 ( .I1(n12668), .I2(n10905), .O(n10754) );
  OA12HHD U8292 ( .B1(n13010), .B2(n7484), .A1(n13458), .O(n7798) );
  ND2HHD U8293 ( .I1(n13478), .I2(n9806), .O(n8794) );
  NR2EHD U8294 ( .I1(n12370), .I2(n12371), .O(n12372) );
  OA13HHD U8295 ( .B1(n10708), .B2(n11467), .B3(n11013), .A1(n12491), .O(n10709) );
  XNR2HHD U8296 ( .I1(n7577), .I2(n9637), .O(n13897) );
  AN3HHD U8297 ( .I1(n10198), .I2(n13058), .I3(n11634), .O(n8213) );
  ND3EHD U8298 ( .I1(n12610), .I2(n11254), .I3(n12640), .O(n11072) );
  NR2CHD U8299 ( .I1(n10587), .I2(n8801), .O(n11181) );
  ND2HHD U8300 ( .I1(n6753), .I2(n9679), .O(n11932) );
  ND3CHD U8301 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(n10562), .I3(n14950), .O(n7620) );
  NR2CHD U8302 ( .I1(n9524), .I2(n9522), .O(n9521) );
  ND3EHD U8303 ( .I1(n9665), .I2(n8900), .I3(n6846), .O(n8568) );
  INVMHD U8304 ( .I(n6714), .O(n7864) );
  ND3EHD U8305 ( .I1(n7016), .I2(n8789), .I3(n8199), .O(n6714) );
  BUFMHD U8306 ( .I(n11022), .O(n9738) );
  BUFNHD U8307 ( .I(n11022), .O(n9897) );
  INVKHD U8308 ( .I(n6905), .O(n10057) );
  INVLHD U8309 ( .I(n10176), .O(n8176) );
  ND2HHD U8310 ( .I1(n6715), .I2(n13827), .O(n9220) );
  NR2GHD U8311 ( .I1(n7939), .I2(n13666), .O(n6715) );
  INVDHD U8312 ( .I(n13926), .O(n7790) );
  INVKHD U8313 ( .I(n6717), .O(n10425) );
  ND2HHD U8314 ( .I1(n12713), .I2(n9723), .O(n6717) );
  NR2GHD U8315 ( .I1(n9911), .I2(n10210), .O(n12357) );
  INVCKGHD U8316 ( .I(n8264), .O(n6718) );
  ND3EHD U8317 ( .I1(n10209), .I2(n8763), .I3(n10107), .O(n6860) );
  NR2IHD U8318 ( .I1(n9947), .I2(n9945), .O(n9864) );
  ND3EHD U8319 ( .I1(n11662), .I2(_i_CLEFIA128_rndcnt_reg _0), .I3(n14927), .O(n11663) );
  INVMHD U8320 ( .I(n7905), .O(n10738) );
  ND2KHD U8321 ( .I1(n6721), .I2(n9844), .O(n7905) );
  BUFEHD U8322 ( .I(n6898), .O(n6722) );
  ND2HHD U8323 ( .I1(n10855), .I2(n6806), .O(n10857) );
  INVNHD U8324 ( .I(_i_CLEFIA128_keyL _74), .O(n8974) );
  INVCKGHD U8325 ( .I(n13550), .O(n7861) );
  ND2KHD U8326 ( .I1(n7930), .I2(n7036), .O(n13550) );
  INVGHD U8327 ( .I(n6887), .O(n8009) );
  ND3EHD U8328 ( .I1(n7490), .I2(n7489), .I3(n7495), .O(n7494) );
  OA13EHD U8329 ( .B1(n12607), .B2(n10852), .B3(n11057), .A1(n11230), .O(n10853) );
  ND2HHD U8330 ( .I1(n8350), .I2(n9146), .O(n12607) );
  ND2KHD U8331 ( .I1(n12497), .I2(n7639), .O(n7209) );
  XNR2KHD U8332 ( .I1(n7640), .I2(n6900), .O(n7639) );
  ND3EHD U8333 ( .I1(n9542), .I2(n12149), .I3(n11735), .O(n11738) );
  INVGHD U8334 ( .I(n12758), .O(n10068) );
  ND3EHD U8335 ( .I1(n12570), .I2(n7278), .I3(n7277), .O(n7276) );
  NR2GHD U8336 ( .I1(n7712), .I2(n7711), .O(n7944) );
  ND2HHD U8337 ( .I1(n8705), .I2(n8312), .O(n8704) );
  ND3CHD U8338 ( .I1(n8704), .I2(n8703), .I3(n14340), .O(n6155) );
  ND3CHD U8339 ( .I1(n14075), .I2(n14074), .I3(n14073), .O(n14077) );
  ND2DHD U8340 ( .I1(n9042), .I2(n10011), .O(n11068) );
  ND2HHD U8341 ( .I1(n7187), .I2(n8202), .O(n11241) );
  NR2GHD U8342 ( .I1(n11242), .I2(n11241), .O(n11243) );
  INVKHD U8343 ( .I(n10446), .O(n9844) );
  ND2KHD U8344 ( .I1(n8914), .I2(n8888), .O(n10731) );
  INVQHD U8345 ( .I(_i_CLEFIA128_keyL _73), .O(n9528) );
  NR2IHD U8346 ( .I1(n9671), .I2(n10077), .O(n7828) );
  BUFEHD U8347 ( .I(n8899), .O(n6724) );
  ND2KHD U8348 ( .I1(n7825), .I2(n7420), .O(n12832) );
  ND2HHD U8349 ( .I1(n10851), .I2(n10850), .O(n8042) );
  ND2KHD U8350 ( .I1(n10794), .I2(n10874), .O(n10850) );
  ND2HHD U8351 ( .I1(n11822), .I2(n11821), .O(n11823) );
  BUFEHD U8352 ( .I(n12511), .O(n6726) );
  ND2HHD U8353 ( .I1(n11510), .I2(n11503), .O(n6728) );
  ND2HHD U8354 ( .I1(n12561), .I2(n9801), .O(n6729) );
  OA12HHD U8355 ( .B1(n7282), .B2(n12557), .A1(n12747), .O(n7281) );
  ND2KHD U8356 ( .I1(n12030), .I2(n13132), .O(n13199) );
  OA12HHD U8357 ( .B1(n15074), .B2(_i_CLEFIA128_keyK _123), .A1(n14405), .O(n11578) );
  AN2HHD U8358 ( .I1(n7187), .I2(n12618), .O(n8444) );
  ND3EHD U8359 ( .I1(n7329), .I2(n10233), .I3(n7328), .O(n7324) );
  INVQHD U8360 ( .I(_i_CLEFIA128_rndcnt_reg _0), .O(n8589) );
  ND3EHD U8361 ( .I1(n7646), .I2(_i_CLEFIA128_rndcnt_reg _0), .I3(_i_CLEFIA128_keyK _35), .O(n7645) );
  ND2HHD U8362 ( .I1(n6730), .I2(_i_CLEFIA128_state_reg _1), .O(n7651) );
  ND3EHD U8363 ( .I1(n7566), .I2(_i_CLEFIA128_rndcnt_reg _0), .I3(n15300), .O(n6730) );
  ND2HHD U8364 ( .I1(n12611), .I2(n12655), .O(n12511) );
  ND2HHD U8365 ( .I1(n10849), .I2(n11250), .O(n8043) );
  ND2KHD U8366 ( .I1(n8791), .I2(n10271), .O(n10849) );
  INVJHD U8367 ( .I(n12496), .O(n11525) );
  INVDHD U8368 ( .I(n10464), .O(n10060) );
  NR2EHD U8369 ( .I1(n8892), .I2(n12052), .O(n8891) );
  INVMHD U8370 ( .I(_i_CLEFIA128_keyL _90), .O(n10031) );
  AN2HHD U8371 ( .I1(n12376), .I2(n12280), .O(n7008) );
  NR2CHD U8372 ( .I1(n8527), .I2(n8804), .O(n7719) );
  ND2HHD U8373 ( .I1(n7522), .I2(n10440), .O(n8804) );
  OAI12CHD U8374 ( .B1(n9979), .B2(n12275), .A1(n13634), .O(n6731) );
  ND2KHD U8375 ( .I1(n9626), .I2(n9087), .O(n12451) );
  OA12HHD U8376 ( .B1(n15069), .B2(_i_CLEFIA128_keyK _81), .A1(n14405), .O(n10564) );
  ND3EHD U8377 ( .I1(n6732), .I2(n7219), .I3(_i_CLEFIA128_rndcnt_reg _0), .O(n8097) );
  ND2HHD U8378 ( .I1(_i_CLEFIA128_keyL _17), .I2(_i_CLEFIA128_keyK _17), .O(n6733) );
  INVGHD U8379 ( .I(n12670), .O(n8594) );
  NR2IHD U8380 ( .I1(n9787), .I2(n9786), .O(n7289) );
  AN3HHD U8381 ( .I1(n13573), .I2(n12401), .I3(n13603), .O(n13153) );
  ND3EHD U8382 ( .I1(n12069), .I2(n11795), .I3(n12298), .O(n11797) );
  ND2DHD U8383 ( .I1(n14053), .I2(n14071), .O(n11622) );
  INVMHD U8384 ( .I(n7200), .O(n6818) );
  OR3HHD U8385 ( .I1(n8073), .I2(n11752), .I3(n11751), .O(n8829) );
  ND2KHD U8386 ( .I1(n13099), .I2(n9631), .O(n11752) );
  OA13EHD U8387 ( .B1(n13675), .B2(n11810), .B3(n13825), .A1(n13817), .O(n7582) );
  ND3EHD U8388 ( .I1(n11800), .I2(n11798), .I3(n11799), .O(n13825) );
  ND2KHD U8389 ( .I1(n9897), .I2(n9898), .O(n11365) );
  NR2GHD U8390 ( .I1(n6738), .I2(n11753), .O(n6737) );
  INVJHD U8391 ( .I(n11821), .O(n6738) );
  INVMHD U8392 ( .I(n7076), .O(n7841) );
  ND2KHD U8393 ( .I1(n7429), .I2(n7050), .O(n7916) );
  NR2IHD U8394 ( .I1(n9036), .I2(n11497), .O(n11498) );
  AN3HHD U8395 ( .I1(n9075), .I2(n9965), .I3(n9967), .O(n6739) );
  XNR2KHD U8396 ( .I1(_i_CLEFIA128_CON_T_xi _9), .I2(DOUT_122), .O(n10188));
  BUFKHD U8397 ( .I(n6899), .O(n6741) );
  AN3B1HHD U8398 ( .I1(n8358), .I2(n13085), .B1(n7334), .O(n8245) );
  ND2KHD U8399 ( .I1(n7915), .I2(n6903), .O(n7015) );
  ND2HHD U8400 ( .I1(n11589), .I2(_i_CLEFIA128_state_reg _1), .O(n8849) );
  ND2KHD U8401 ( .I1(n9438), .I2(n9437), .O(n9404) );
  ND2KHD U8402 ( .I1(n9832), .I2(n8866), .O(n12108) );
  BUFKHD U8403 ( .I(n7965), .O(n6742) );
  NR2IHD U8404 ( .I1(n9214), .I2(n12975), .O(n11907) );
  ND3EHD U8405 ( .I1(n6743), .I2(n9227), .I3(n9228), .O(n9226) );
  ND3EHD U8406 ( .I1(n11757), .I2(n11756), .I3(n13241), .O(n6743) );
  ND2HHD U8407 ( .I1(n8367), .I2(n6744), .O(n10559) );
  INVCKGHD U8408 ( .I(n8798), .O(n6745) );
  ND2KHD U8409 ( .I1(n9087), .I2(n9017), .O(n10978) );
  ND2KHD U8410 ( .I1(n6746), .I2(n7677), .O(n9700) );
  NR2IHD U8411 ( .I1(n7014), .I2(n7674), .O(n6746) );
  ND2KHD U8412 ( .I1(n13837), .I2(n9210), .O(n11706) );
  ND2KHD U8413 ( .I1(n12423), .I2(n12327), .O(n13365) );
  OR2B1CHD U8414 ( .I1(_i_CLEFIA128_keyK _63), .B1(n10337), .O(n11596) );
  ND3EHD U8415 ( .I1(n6749), .I2(n6747), .I3(n8131), .O(n11600) );
  ND2HHD U8416 ( .I1(n11598), .I2(n6748), .O(n6747) );
  ND2HHD U8417 ( .I1(n11597), .I2(_i_CLEFIA128_keyL _63), .O(n6749) );
  ND3EHD U8418 ( .I1(n8826), .I2(n10308), .I3(n10309), .O(n7852) );
  ND2HHD U8419 ( .I1(n7580), .I2(n7606), .O(n12529) );
  AN2EHD U8420 ( .I1(n12610), .I2(n12611), .O(n6792) );
  NR2GHD U8421 ( .I1(n6751), .I2(n6750), .O(n8237) );
  ND3EHD U8422 ( .I1(n12497), .I2(n7639), .I3(n8801), .O(n6751) );
  ND3EHD U8423 ( .I1(n6752), .I2(n7634), .I3(n7636), .O(n12373) );
  ND3EHD U8424 ( .I1(n7633), .I2(n12349), .I3(n7632), .O(n6752) );
  BUFKHD U8425 ( .I(n12366), .O(n6753) );
  ND2KHD U8426 ( .I1(n7104), .I2(n10687), .O(n14137) );
  OA22HHD U8427 ( .A1(n10686), .A2(n10685), .B1(n10684), .B2(n10683), .O(n7104) );
  ND2HHD U8428 ( .I1(n8656), .I2(n9886), .O(n12110) );
  BUFHHD U8429 ( .I(n12914), .O(n8897) );
  AN2HHD U8430 ( .I1(n11235), .I2(n9648), .O(n6812) );
  OR3HHD U8431 ( .I1(n10865), .I2(n10863), .I3(n10864), .O(n10866) );
  NR2GHD U8432 ( .I1(n8954), .I2(n6754), .O(n7768) );
  ND2HHD U8433 ( .I1(n12842), .I2(n6917), .O(n6754) );
  ND2KHD U8434 ( .I1(n15281), .I2(_i_CLEFIA128_rndcnt_reg _0), .O(n6844) );
  ND2HHD U8435 ( .I1(n10971), .I2(n6716), .O(n8542) );
  NR3BHD U8436 ( .I1(n11432), .I2(n7913), .I3(n11461), .O(n6853) );
  ND3EHD U8437 ( .I1(n8161), .I2(n8872), .I3(n11988), .O(n8160) );
  XOR2HHD U8438 ( .I1(n10455), .I2(n6756), .O(n9802) );
  ND2HHD U8439 ( .I1(n7087), .I2(n7086), .O(n6756) );
  NR2IHD U8440 ( .I1(n6757), .I2(n7892), .O(n10240) );
  ND2KHD U8441 ( .I1(n9218), .I2(n11530), .O(n6757) );
  ND3EHD U8442 ( .I1(n9789), .I2(_i_CLEFIA128_rndcnt_reg _0), .I3(n15257), .O(n8745) );
  ND2KHD U8443 ( .I1(_i_CLEFIA128_keyK _5), .I2(n8797), .O(n9789) );
  ND2KHD U8444 ( .I1(n7219), .I2(_i_CLEFIA128_keyK _24), .O(n9418) );
  INVQHD U8445 ( .I(n8798), .O(n7219) );
  ND3EHD U8446 ( .I1(n8544), .I2(n8543), .I3(n14166), .O(n6194) );
  ND3EHD U8447 ( .I1(n7995), .I2(n8802), .I3(n8857), .O(n7994) );
  ND2HHD U8448 ( .I1(n6758), .I2(n10060), .O(n10059) );
  ND2HHD U8449 ( .I1(n10243), .I2(n10244), .O(n6758) );
  XNR2HHD U8450 ( .I1(n9442), .I2(n7479), .O(n10176) );
  ND2KHD U8451 ( .I1(n7481), .I2(n7480), .O(n7479) );
  BUFMHD U8452 ( .I(n12373), .O(n14329) );
  NR2GHD U8453 ( .I1(n7295), .I2(n7296), .O(n10146) );
  OA13EHD U8454 ( .B1(n11293), .B2(n12508), .B3(n12492), .A1(n12474), .O(n11294) );
  NR2GHD U8455 ( .I1(n10445), .I2(n7783), .O(n10293) );
  ND2HHD U8456 ( .I1(n8504), .I2(n8499), .O(n8896) );
  ND2HHD U8457 ( .I1(n11887), .I2(_i_CLEFIA128_state_reg _1), .O(n6759) );
  NR2IHD U8458 ( .I1(n10431), .I2(n7338), .O(n7337) );
  ND2KHD U8459 ( .I1(n10441), .I2(n10767), .O(n7338) );
  OA13EHD U8460 ( .B1(n12515), .B2(n12514), .B3(n7485), .A1(n12662), .O(n12551) );
  ND3EHD U8461 ( .I1(n9378), .I2(n6761), .I3(n6760), .O(n8723) );
  INVGHD U8462 ( .I(n10758), .O(n6761) );
  ND2HHD U8463 ( .I1(n8657), .I2(n13582), .O(n8706) );
  OR2KHD U8464 ( .I1(n8801), .I2(n7990), .O(n8211) );
  ND2HHD U8465 ( .I1(n10281), .I2(n10583), .O(n7990) );
  XNR2HHD U8466 ( .I1(DOUT_4), .I2(n14137), .O(n8517) );
  INVKHD U8467 ( .I(n10474), .O(n7133) );
  ND2KHD U8468 ( .I1(n6819), .I2(n12749), .O(n7664) );
  ND3EHD U8469 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(n7069), .I3(n14954), .O(n8702) );
  MUX2HHD U8470 ( .A(n13885), .B(n13884), .S(n15439), .O(n8805) );
  XNR2KHD U8471 ( .I1(n13883), .I2(n6762), .O(n15439) );
  XOR2HHD U8472 ( .I1(n8806), .I2(n14493), .O(n6762) );
  INVKHD U8473 ( .I(n6763), .O(n8233) );
  ND3EHD U8474 ( .I1(n8508), .I2(n8977), .I3(n8547), .O(n6763) );
  NR2IHD U8475 ( .I1(n8798), .I2(n7575), .O(n7576) );
  XNR2KHD U8476 ( .I1(_i_CLEFIA128_keyL _65), .I2(n8001), .O(n10465) );
  OA112EHD U8477 ( .C1(n11877), .C2(n8679), .A1(n8678), .B1(_i_CLEFIA128_state_reg _1), .O(n8677) );
  BUFKHD U8478 ( .I(n9359), .O(n6764) );
  BUFEHD U8479 ( .I(n7042), .O(n6766) );
  ND2KHD U8480 ( .I1(n8938), .I2(n10219), .O(n10818) );
  BUFEHD U8481 ( .I(n10761), .O(n6767) );
  OR3HHD U8482 ( .I1(n13243), .I2(n13225), .I3(n13224), .O(n13226) );
  NR2CHD U8483 ( .I1(n10643), .I2(n6768), .O(n9711) );
  ND3EHD U8484 ( .I1(n6769), .I2(n9713), .I3(n12513), .O(n6768) );
  INVGHD U8485 ( .I(n10642), .O(n6769) );
  BUFKHD U8486 ( .I(n9678), .O(n6770) );
  ND2HHD U8487 ( .I1(n7222), .I2(n6972), .O(n10951) );
  NR2GHD U8488 ( .I1(n10136), .I2(n10137), .O(n11204) );
  NR2GHD U8489 ( .I1(n11205), .I2(n10801), .O(n9618) );
  ND2KHD U8490 ( .I1(n7859), .I2(n13643), .O(n7929) );
  ND2HHD U8491 ( .I1(n8798), .I2(_i_CLEFIA128_keyL _68), .O(n10459) );
  XNR2KHD U8492 ( .I1(n8651), .I2(n13973), .O(n8553) );
  OR2EHD U8493 ( .I1(n6776), .I2(n10339), .O(n6775) );
  ND2HHD U8494 ( .I1(n7350), .I2(n7351), .O(n6777) );
  INVCKIHD U8495 ( .I(n8425), .O(n9924) );
  ND2KHD U8496 ( .I1(n9807), .I2(n7933), .O(n13842) );
  ND2HHD U8497 ( .I1(n7374), .I2(n7184), .O(n9997) );
  ND2HHD U8498 ( .I1(n11990), .I2(n7389), .O(n10113) );
  NR2GHD U8499 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(n6779), .O(n9091) );
  ND2HHD U8500 ( .I1(n9752), .I2(n9126), .O(n12113) );
  ND2HHD U8501 ( .I1(n8511), .I2(n10759), .O(n8813) );
  ND2DHD U8502 ( .I1(n9113), .I2(n6780), .O(n9112) );
  NR3BHD U8503 ( .I1(n13465), .I2(n13464), .I3(n13466), .O(n6780) );
  NR2EHD U8504 ( .I1(n12099), .I2(n12098), .O(n12100) );
  NR2IHD U8505 ( .I1(n7546), .I2(n7361), .O(n11090) );
  NR2EHD U8506 ( .I1(n12851), .I2(n10826), .O(n10832) );
  ND2HHD U8507 ( .I1(n8466), .I2(n8450), .O(n8465) );
  ND2DHD U8508 ( .I1(n8607), .I2(n8018), .O(n11393) );
  ND3EHD U8509 ( .I1(n9334), .I2(n13429), .I3(n9338), .O(n7140) );
  ND3EHD U8510 ( .I1(n6781), .I2(n7317), .I3(n12605), .O(n10639) );
  INVGHD U8511 ( .I(n6782), .O(n6781) );
  ND3CHD U8512 ( .I1(n11262), .I2(n11063), .I3(n10850), .O(n6782) );
  ND2DHD U8513 ( .I1(n13222), .I2(n8061), .O(n13105) );
  ND2DHD U8514 ( .I1(n10001), .I2(n8217), .O(n6200) );
  XOR2HHD U8515 ( .I1(_i_CLEFIA128_keyL _109), .I2(n11889), .O(n11891) );
  INVNHD U8516 ( .I(n9102), .O(n8209) );
  NR2GHD U8517 ( .I1(n12761), .I2(n6783), .O(n6849) );
  ND3EHD U8518 ( .I1(n9094), .I2(n6677), .I3(n13680), .O(n13683) );
  ND2HHD U8519 ( .I1(n9847), .I2(n13398), .O(n12421) );
  INVKHD U8520 ( .I(n11905), .O(n8126) );
  AN3HHD U8521 ( .I1(n11529), .I2(n12486), .I3(n9531), .O(n7004) );
  INVJHD U8522 ( .I(n12185), .O(n9646) );
  NR2GHD U8523 ( .I1(n9671), .I2(n11072), .O(n12604) );
  AN3B1HHD U8524 ( .I1(n6894), .I2(n9034), .B1(n6784), .O(n11418) );
  INVKHD U8525 ( .I(n11811), .O(n7641) );
  ND2HHD U8526 ( .I1(n10794), .I2(n9766), .O(n10862) );
  NR2GHD U8527 ( .I1(n12308), .I2(n12307), .O(n12311) );
  OR3HHD U8528 ( .I1(n12758), .I2(n12757), .I3(n12756), .O(n12760) );
  INVQHD U8529 ( .I(n7991), .O(n9050) );
  AN2HHD U8530 ( .I1(n7967), .I2(n8253), .O(n6934) );
  BUFGHD U8531 ( .I(n11504), .O(n7099) );
  ND3CHD U8532 ( .I1(n9726), .I2(n12220), .I3(n13365), .O(n12221) );
  XNR2KHD U8533 ( .I1(n6786), .I2(n6787), .O(n9817) );
  XOR2EHD U8534 ( .I1(DOUT_85), .I2(n9519), .O(n6786) );
  NR2IHD U8535 ( .I1(n9555), .I2(n9554), .O(n10239) );
  ND2KHD U8536 ( .I1(n10619), .I2(n7053), .O(n8775) );
  AN2HHD U8537 ( .I1(n12621), .I2(n10847), .O(n10837) );
  OR3CHD U8538 ( .I1(n13481), .I2(n7764), .I3(n13480), .O(n13485) );
  AN2HHD U8539 ( .I1(n11592), .I2(n6796), .O(n8355) );
  ND2HHD U8540 ( .I1(n10215), .I2(n9539), .O(n6788) );
  ND2HHD U8541 ( .I1(n6535), .I2(n6897), .O(n12034) );
  ND2KHD U8542 ( .I1(n12902), .I2(n10095), .O(n6897) );
  ND2HHD U8543 ( .I1(n11271), .I2(n11270), .O(n8486) );
  BUFGHD U8544 ( .I(n11547), .O(n9591) );
  AN2HHD U8545 ( .I1(n11814), .I2(n13804), .O(n6960) );
  ND3CHD U8546 ( .I1(n13088), .I2(n13085), .I3(n8197), .O(n11652) );
  NR2IHD U8547 ( .I1(n7889), .I2(n10967), .O(n7888) );
  NR2EHD U8548 ( .I1(n10957), .I2(n10967), .O(n10753) );
  ND2KHD U8549 ( .I1(n10152), .I2(n7783), .O(n9327) );
  ND2DHD U8550 ( .I1(n8337), .I2(n12790), .O(n7476) );
  AN3HHD U8551 ( .I1(n8194), .I2(n8337), .I3(n10899), .O(n12705) );
  AN2B1CHD U8552 ( .I1(n8337), .B1(n12809), .O(n12810) );
  ND2KHD U8553 ( .I1(n9559), .I2(n7420), .O(n8337) );
  ND2HHD U8554 ( .I1(n11766), .I2(n7335), .O(n11644) );
  AN2EHD U8555 ( .I1(n10619), .I2(n8179), .O(n6929) );
  ND2HHD U8556 ( .I1(n11834), .I2(n11763), .O(n9556) );
  INVMHD U8557 ( .I(n9918), .O(n9458) );
  ND3EHD U8558 ( .I1(n8442), .I2(n6587), .I3(n14070), .O(n11657) );
  ND2HHD U8559 ( .I1(n12612), .I2(n6792), .O(n12613) );
  BUFLHD U8560 ( .I(n11548), .O(n9733) );
  ND2HHD U8561 ( .I1(n9738), .I2(n11095), .O(n12736) );
  NR2EHD U8562 ( .I1(n11084), .I2(n11085), .O(n11086) );
  ND3EHD U8563 ( .I1(n6793), .I2(n6795), .I3(n6794), .O(n7126) );
  AN3EHD U8564 ( .I1(n10511), .I2(n11376), .I3(n10510), .O(n6794) );
  NR3BHD U8565 ( .I1(n12721), .I2(n12720), .I3(n11038), .O(n6795) );
  INVNHD U8566 ( .I(n11647), .O(n13058) );
  AN2EHD U8567 ( .I1(n7394), .I2(n11647), .O(n8027) );
  INVMHD U8568 ( .I(n7721), .O(n8133) );
  NR2IHD U8569 ( .I1(n10479), .I2(n12748), .O(n10480) );
  AN2EHD U8570 ( .I1(n12558), .I2(n11323), .O(n10507) );
  INVNHD U8571 ( .I(n8589), .O(n9173) );
  ND2DHD U8572 ( .I1(n9423), .I2(n12622), .O(n10871) );
  AN2HHD U8573 ( .I1(n10441), .I2(n10431), .O(n8397) );
  NR2EHD U8574 ( .I1(n11265), .I2(n10014), .O(n11266) );
  NR2GHD U8575 ( .I1(n8804), .I2(n8501), .O(n8500) );
  ND2DHD U8576 ( .I1(n10813), .I2(n10810), .O(n8503) );
  ND3CHD U8577 ( .I1(n12566), .I2(n8101), .I3(n7309), .O(n12567) );
  ND2KHD U8578 ( .I1(n11142), .I2(n6893), .O(n9765) );
  OR3EHD U8579 ( .I1(n11422), .I2(n11421), .I3(n11420), .O(n11428) );
  NR2GHD U8580 ( .I1(n11154), .I2(n9045), .O(n11200) );
  NR2GHD U8581 ( .I1(n7863), .I2(n10328), .O(n10791) );
  INVKHD U8582 ( .I(n12189), .O(n7093) );
  ND3EHD U8583 ( .I1(n8983), .I2(n6993), .I3(n8344), .O(n6797) );
  XOR2HHD U8584 ( .I1(n8561), .I2(n13972), .O(n6798) );
  ND2DHD U8585 ( .I1(n8515), .I2(n11485), .O(n11391) );
  NR2IHD U8586 ( .I1(n11280), .I2(n10594), .O(n10598) );
  ND2DHD U8587 ( .I1(n7704), .I2(n8078), .O(n14042) );
  AN2HHD U8588 ( .I1(n11967), .I2(n9884), .O(n6799) );
  ND2HHD U8589 ( .I1(n8710), .I2(n13622), .O(n8709) );
  ND2KHD U8590 ( .I1(n11628), .I2(n11840), .O(n9493) );
  INVGHD U8591 ( .I(n11265), .O(n11261) );
  INVQHD U8592 ( .I(n7477), .O(n10179) );
  NR2EHD U8593 ( .I1(n9337), .I2(n9336), .O(n9335) );
  ND3EHD U8594 ( .I1(n8266), .I2(n13439), .I3(n6986), .O(n9336) );
  XNR3EHD U8595 ( .I1(n13741), .I2(n9797), .I3(n6800), .O(n6802) );
  AN2HHD U8596 ( .I1(n9694), .I2(n8014), .O(n6951) );
  ND2HHD U8597 ( .I1(n6895), .I2(n9694), .O(n12581) );
  AN2EHD U8598 ( .I1(n7897), .I2(n9568), .O(n6801) );
  NR2EHD U8599 ( .I1(n9055), .I2(n11066), .O(n9054) );
  ND2KHD U8600 ( .I1(n8896), .I2(n9849), .O(n13951) );
  XOR2HHD U8601 ( .I1(n13266), .I2(n6802), .O(n8067) );
  OA112EHD U8602 ( .C1(n6875), .C2(n13218), .A1(n13066), .B1(n14071), .O(n13071) );
  AN3EHD U8603 ( .I1(n14071), .I2(n6641), .I3(n7077), .O(n14054) );
  INVMHD U8604 ( .I(n10587), .O(n10583) );
  INVKHD U8605 ( .I(n11775), .O(n7041) );
  NR2IHD U8606 ( .I1(n12627), .I2(n10646), .O(n12513) );
  ND3CHD U8607 ( .I1(n7365), .I2(n12662), .I3(n6841), .O(n10643) );
  BUFNHD U8608 ( .I(n10111), .O(n7671) );
  XOR2KHD U8609 ( .I1(n10343), .I2(n10342), .O(n6803) );
  NR2GHD U8610 ( .I1(n12151), .I2(n12152), .O(n12321) );
  NR2EHD U8611 ( .I1(n12151), .I2(n12143), .O(n11780) );
  NR2IHD U8612 ( .I1(n11294), .I2(n9052), .O(n9782) );
  INVKHD U8613 ( .I(n13098), .O(n13244) );
  INVGHD U8614 ( .I(n10850), .O(n11224) );
  ND2DHD U8615 ( .I1(n15171), .I2(n11130), .O(n9107) );
  NR2IHD U8616 ( .I1(n10474), .I2(n7132), .O(n12750) );
  INVNHD U8617 ( .I(n6804), .O(n6805) );
  NR2GHD U8618 ( .I1(n12700), .I2(n12699), .O(n12863) );
  ND2HHD U8619 ( .I1(n12030), .I2(n12383), .O(n13134) );
  AN2EHD U8620 ( .I1(n12030), .I2(n7648), .O(n12279) );
  ND2DHD U8621 ( .I1(n8914), .I2(n12692), .O(n12693) );
  NR2EHD U8622 ( .I1(n12694), .I2(n12693), .O(n12697) );
  NR2GHD U8623 ( .I1(n11547), .I2(n11166), .O(n10111) );
  ND2HHD U8624 ( .I1(n11522), .I2(n11440), .O(n11177) );
  ND2KHD U8625 ( .I1(n6562), .I2(n11948), .O(n9693) );
  INVCKIHD U8626 ( .I(n13241), .O(n11640) );
  ND2HHD U8627 ( .I1(n14076), .I2(n13222), .O(n8128) );
  ND2HHD U8628 ( .I1(n13383), .I2(n13036), .O(n11956) );
  INVDHD U8629 ( .I(n8188), .O(n7498) );
  OA112HHD U8630 ( .C1(n6899), .C2(n11868), .A1(n11867), .B1(_i_CLEFIA128_state_reg _1), .O(n11872) );
  OR2EHD U8631 ( .I1(n10358), .I2(n9997), .O(n8334) );
  ND3EHD U8632 ( .I1(n10711), .I2(n10988), .I3(n11534), .O(n10985) );
  NR2EHD U8633 ( .I1(n8094), .I2(n7026), .O(n10711) );
  BUFQHD U8634 ( .I(n11897), .O(n12251) );
  NR2IHD U8635 ( .I1(n7182), .I2(n10383), .O(n7122) );
  AN3EHD U8636 ( .I1(n7206), .I2(n11411), .I3(n11340), .O(n10518) );
  NR2GHD U8637 ( .I1(n10743), .I2(n9382), .O(n9381) );
  NR2IHD U8638 ( .I1(n10709), .I2(n10726), .O(n9935) );
  ND3HHD U8639 ( .I1(n10971), .I2(n8564), .I3(n6716), .O(n8365) );
  INVDHD U8640 ( .I(n10902), .O(n8814) );
  AN3HHD U8641 ( .I1(n9111), .I2(n7003), .I3(n7002), .O(n6807) );
  INVNHD U8642 ( .I(n7334), .O(n13478) );
  NR2EHD U8643 ( .I1(n11144), .I2(n11143), .O(n11145) );
  ND2KHD U8644 ( .I1(n10096), .I2(n8286), .O(n9018) );
  ND3EHD U8645 ( .I1(n12114), .I2(n12284), .I3(n12948), .O(n12115) );
  ND3EHD U8646 ( .I1(n7668), .I2(n12776), .I3(n10053), .O(n7667) );
  ND2KHD U8647 ( .I1(n7161), .I2(n10668), .O(n10851) );
  INVDHD U8648 ( .I(n12493), .O(n8822) );
  INVKHD U8649 ( .I(n9582), .O(n11183) );
  ND3EHD U8650 ( .I1(n11291), .I2(n12473), .I3(n11290), .O(n11293) );
  INVJHD U8651 ( .I(n12598), .O(n11073) );
  NR2GHD U8652 ( .I1(n6931), .I2(n10051), .O(n10037) );
  ND2DHD U8653 ( .I1(n7417), .I2(n13592), .O(n7468) );
  ND2HHD U8654 ( .I1(n7417), .I2(n13130), .O(n7550) );
  ND2HHD U8655 ( .I1(n12788), .I2(n8547), .O(n9361) );
  ND2HHD U8656 ( .I1(n6893), .I2(n9116), .O(n10585) );
  ND2HHD U8657 ( .I1(n8226), .I2(n9455), .O(n12208) );
  OA12EHD U8658 ( .B1(n7524), .B2(n12840), .A1(n7523), .O(n6809) );
  NR2EHD U8659 ( .I1(n13061), .I2(n13224), .O(n13063) );
  ND2DHD U8660 ( .I1(n12794), .I2(n9559), .O(n12710) );
  ND2HHD U8661 ( .I1(n10739), .I2(n9559), .O(n12878) );
  NR2EHD U8662 ( .I1(n10869), .I2(n10792), .O(n10800) );
  ND3EHD U8663 ( .I1(n13371), .I2(n12427), .I3(n12426), .O(n12429) );
  ND3CHD U8664 ( .I1(n12570), .I2(n12763), .I3(n11377), .O(n11388) );
  NR2EHD U8665 ( .I1(n11469), .I2(n9086), .O(n11354) );
  ND2HHD U8666 ( .I1(n13102), .I2(n8061), .O(n8060) );
  ND2HHD U8667 ( .I1(n12646), .I2(n6812), .O(n10679) );
  ND2HHD U8668 ( .I1(n6883), .I2(n10773), .O(n11235) );
  ND2KHD U8669 ( .I1(n9287), .I2(n12462), .O(n9967) );
  AN2HHD U8670 ( .I1(n11216), .I2(n11245), .O(n12662) );
  ND2KHD U8671 ( .I1(n13078), .I2(n9631), .O(n12195) );
  ND3EHD U8672 ( .I1(n13078), .I2(n13469), .I3(n14067), .O(n8598) );
  ND2HHD U8673 ( .I1(n13078), .I2(n13470), .O(n7716) );
  ND3CHD U8674 ( .I1(n13098), .I2(n14082), .I3(n14083), .O(n13061) );
  ND2DHD U8675 ( .I1(n11443), .I2(n12454), .O(n11444) );
  AN2HHD U8676 ( .I1(n12454), .I2(n12453), .O(n12455) );
  AN3EHD U8677 ( .I1(n12454), .I2(n9359), .I3(n11191), .O(n10722) );
  BUFGHD U8678 ( .I(n7488), .O(n7199) );
  ND2HHD U8679 ( .I1(n7580), .I2(n11062), .O(n10634) );
  INVKHD U8680 ( .I(n10425), .O(n7747) );
  ND2HHD U8681 ( .I1(n12562), .I2(n8188), .O(n8452) );
  ND2HHD U8682 ( .I1(n11155), .I2(n9144), .O(n10595) );
  ND2HHD U8683 ( .I1(n10891), .I2(n7730), .O(n7729) );
  ND2KHD U8684 ( .I1(n9066), .I2(n9105), .O(n6816) );
  ND2HHD U8685 ( .I1(n9066), .I2(n9105), .O(n14170) );
  ND2HHD U8686 ( .I1(n8183), .I2(n11995), .O(n12920) );
  BUFQHD U8687 ( .I(n7474), .O(n7420) );
  NR2IHD U8688 ( .I1(n9568), .I2(n7500), .O(n9422) );
  AN2EHD U8689 ( .I1(n8232), .I2(n10966), .O(n10881) );
  XNR2KHD U8690 ( .I1(n14767), .I2(n7505), .O(n7831) );
  NR2IHD U8691 ( .I1(n11074), .I2(n11073), .O(n11217) );
  ND3EHD U8692 ( .I1(n12640), .I2(n11226), .I3(n11068), .O(n9426) );
  NR2GHD U8693 ( .I1(n10735), .I2(n10736), .O(n9638) );
  NR2GHD U8694 ( .I1(n10589), .I2(n10590), .O(n10591) );
  ND2HHD U8695 ( .I1(n8116), .I2(n9050), .O(n6817) );
  ND2HHD U8696 ( .I1(n7621), .I2(n9087), .O(n11541) );
  ND3EHD U8697 ( .I1(n13643), .I2(n12298), .I3(n13550), .O(n11711) );
  AN2B1HHD U8698 ( .I1(n9131), .B1(_i_CLEFIA128_rndcnt_reg _0), .O(n7380) );
  AN2HHD U8699 ( .I1(n8303), .I2(n10885), .O(n8231) );
  ND2KHD U8700 ( .I1(n7474), .I2(n12830), .O(n10959) );
  INVKHD U8701 ( .I(n7596), .O(n12830) );
  NR2IHD U8702 ( .I1(n11928), .I2(n12975), .O(n11898) );
  INVQHD U8703 ( .I(n11911), .O(n12975) );
  ND2HHD U8704 ( .I1(n10858), .I2(n10859), .O(n10860) );
  OA12HHD U8705 ( .B1(n12608), .B2(n9063), .A1(n12605), .O(n9307) );
  ND2DHD U8706 ( .I1(n14066), .I2(n14065), .O(n9400) );
  NR2GHD U8707 ( .I1(n10844), .I2(n10843), .O(n10845) );
  INVJHD U8708 ( .I(n14071), .O(n7290) );
  ND2KHD U8709 ( .I1(n7499), .I2(n12736), .O(n7680) );
  NR2IHD U8710 ( .I1(n7286), .I2(n7274), .O(n13715) );
  AN2HHD U8711 ( .I1(n10329), .I2(n11226), .O(n8431) );
  XNR2HHD U8712 ( .I1(n13953), .I2(n14013), .O(n9962) );
  XOR2KHD U8713 ( .I1(n6788), .I2(n13911), .O(n14804) );
  NR2GHD U8714 ( .I1(n11000), .I2(n9289), .O(n9288) );
  ND2KHD U8715 ( .I1(n7657), .I2(n11491), .O(n11470) );
  ND2HHD U8716 ( .I1(n8245), .I2(n13229), .O(n13230) );
  INVGHD U8717 ( .I(n10017), .O(n10018) );
  XOR3EHD U8718 ( .I1(DOUT_69), .I2(n14215), .I3(n7231), .O(n6821) );
  ND2HHD U8719 ( .I1(n9840), .I2(n7718), .O(n7497) );
  ND2HHD U8720 ( .I1(n11358), .I2(n11349), .O(n11469) );
  INVMHD U8721 ( .I(n12264), .O(n12120) );
  INVKHD U8722 ( .I(n10415), .O(n6822) );
  BUFKHD U8723 ( .I(n9959), .O(n9550) );
  INVMHD U8724 ( .I(n7044), .O(n6823) );
  INVNHD U8725 ( .I(n13058), .O(n7044) );
  XNR2HHD U8726 ( .I1(n8774), .I2(n14489), .O(n8766) );
  ND2HHD U8727 ( .I1(n7791), .I2(n6851), .O(n9448) );
  OR3HHD U8728 ( .I1(n12757), .I2(n11328), .I3(n11327), .O(n11329) );
  INVLHD U8729 ( .I(n8076), .O(n11634) );
  INVGHD U8730 ( .I(n11281), .O(n6854) );
  NR2EHD U8731 ( .I1(n13237), .I2(n13238), .O(n13239) );
  ND2HHD U8732 ( .I1(n9517), .I2(n6742), .O(n13476) );
  NR2IHD U8733 ( .I1(n9367), .I2(n11627), .O(n9517) );
  ND3CHD U8734 ( .I1(n12204), .I2(n14048), .I3(n14074), .O(n8059) );
  OR3HHD U8735 ( .I1(n13488), .I2(n8993), .I3(n13480), .O(n12212) );
  ND2DHD U8736 ( .I1(n8799), .I2(n7384), .O(n9809) );
  INVCHD U8737 ( .I(n12119), .O(n7460) );
  OAI12EHD U8738 ( .B1(n12901), .B2(n12129), .A1(n12125), .O(n12126) );
  ND2KHD U8739 ( .I1(n9020), .I2(n9844), .O(n7230) );
  NR2GHD U8740 ( .I1(n12614), .I2(n12613), .O(n12616) );
  ND3CHD U8741 ( .I1(n7580), .I2(n12621), .I3(n11069), .O(n9005) );
  ND3CHD U8742 ( .I1(n11063), .I2(n12538), .I3(n10778), .O(n10779) );
  ND2DHD U8743 ( .I1(n11063), .I2(n12637), .O(n7193) );
  INVQHD U8744 ( .I(n7316), .O(n10178) );
  AN2HHD U8745 ( .I1(n10415), .I2(n10417), .O(n10201) );
  INVNHD U8746 ( .I(n10281), .O(n9129) );
  XOR2HHD U8747 ( .I1(n9957), .I2(n8651), .O(n9717) );
  ND3CHD U8748 ( .I1(n15404), .I2(n8797), .I3(_i_CLEFIA128_keyK _99), .O(n9884) );
  OA12HHD U8749 ( .B1(n14601), .B2(n15450), .A1(n12897), .O(n10040) );
  ND2KHD U8750 ( .I1(n7389), .I2(n8797), .O(n8130) );
  ND3CHD U8751 ( .I1(n13487), .I2(n13469), .I3(n8061), .O(n11767) );
  ND2HHD U8752 ( .I1(n13470), .I2(n8061), .O(n13080) );
  ND3CHD U8753 ( .I1(n13469), .I2(n8197), .I3(n14043), .O(n7423) );
  OA22HHD U8754 ( .A1(n7924), .A2(n7927), .B1(DOUT_84), .B2(n14342), .O(n9611) );
  INVMHD U8755 ( .I(n9810), .O(n7036) );
  ND2KHD U8756 ( .I1(n7219), .I2(_i_CLEFIA128_keyK _53), .O(n11662) );
  ND2KHD U8757 ( .I1(n7922), .I2(n7923), .O(n9156) );
  ND2DHD U8758 ( .I1(n11296), .I2(n11284), .O(n11140) );
  ND2DHD U8759 ( .I1(n11531), .I2(n11440), .O(n9689) );
  ND2DHD U8760 ( .I1(n9298), .I2(n12487), .O(n7912) );
  ND2DHD U8761 ( .I1(n7376), .I2(n11429), .O(n10996) );
  AN3EHD U8762 ( .I1(n7900), .I2(n11429), .I3(n7304), .O(n7003) );
  ND2HHD U8763 ( .I1(n10945), .I2(n9190), .O(n10901) );
  ND2HHD U8764 ( .I1(n10347), .I2(n6843), .O(n10349) );
  ND3CHD U8765 ( .I1(n10798), .I2(n8202), .I3(n6806), .O(n10650) );
  INVCKIHD U8766 ( .I(n10721), .O(n10593) );
  AN3HHD U8767 ( .I1(n11292), .I2(n12479), .I3(n9224), .O(n10991) );
  ND3EHD U8768 ( .I1(n10753), .I2(n10752), .I3(n10751), .O(n10758) );
  BUFNHD U8769 ( .I(n11707), .O(n9549) );
  AN2KHD U8770 ( .I1(n12053), .I2(n12063), .O(n13608) );
  ND2HHD U8771 ( .I1(n12902), .I2(n12030), .O(n12376) );
  NR2IHD U8772 ( .I1(n7796), .I2(n7795), .O(n7794) );
  XOR2HHD U8773 ( .I1(n8796), .I2(n7363), .O(n14352) );
  INVJHD U8774 ( .I(n8800), .O(n6840) );
  INVDHD U8775 ( .I(n7695), .O(n7687) );
  INVKHD U8776 ( .I(n9821), .O(n9822) );
  ND2DHD U8777 ( .I1(n12469), .I2(n11541), .O(n6826) );
  ND2HHD U8778 ( .I1(n11542), .I2(n6827), .O(n11543) );
  INVDHD U8779 ( .I(n6826), .O(n6827) );
  INVGHD U8780 ( .I(n11420), .O(n11542) );
  NR2GHD U8781 ( .I1(n8599), .I2(n8598), .O(n8597) );
  ND2HHD U8782 ( .I1(n11596), .I2(n6843), .O(n11598) );
  ND2HHD U8783 ( .I1(n15340), .I2(_i_CLEFIA128_rndcnt_reg _0), .O(n6828) );
  ND2HHD U8784 ( .I1(n11570), .I2(n6829), .O(n11571) );
  INVQHD U8785 ( .I(_i_CLEFIA128_keyL _58), .O(n15340) );
  ND2HHD U8786 ( .I1(n11965), .I2(n6796), .O(n11966) );
  XNR2KHD U8787 ( .I1(n6830), .I2(n10418), .O(n8572) );
  ND3EHD U8788 ( .I1(n11526), .I2(n7986), .I3(n6858), .O(n11527) );
  INVQHD U8789 ( .I(_i_CLEFIA128_keyL _75), .O(n6830) );
  ND2HHD U8790 ( .I1(n12714), .I2(n10728), .O(n7732) );
  ND2KHD U8791 ( .I1(n10760), .I2(n7723), .O(n10728) );
  NR2GHD U8792 ( .I1(n9799), .I2(n9161), .O(n9022) );
  OA13EHD U8793 ( .B1(n11468), .B2(n11466), .B3(n11467), .A1(n12462), .O(n9799) );
  OAI12HHD U8794 ( .B1(n9855), .B2(n7420), .A1(n7597), .O(n8425) );
  ND2HHD U8795 ( .I1(n11529), .I2(n9218), .O(n9048) );
  NR2GHD U8796 ( .I1(n12353), .I2(n7442), .O(n7123) );
  NR2IHD U8797 ( .I1(n11928), .I2(n11911), .O(n9450) );
  NR2CHD U8798 ( .I1(n7990), .I2(n7209), .O(n7208) );
  INVCKLHD U8799 ( .I(n14140), .O(n9797) );
  ND2DHD U8800 ( .I1(n14081), .I2(n13076), .O(n13082) );
  ND2HHD U8801 ( .I1(n8797), .I2(_i_CLEFIA128_keyK _36), .O(n11962) );
  BUFKHD U8802 ( .I(n9836), .O(n9779) );
  NR2IHD U8803 ( .I1(n9390), .I2(n9391), .O(n8699) );
  INVGHD U8804 ( .I(n9759), .O(n8623) );
  ND2HHD U8805 ( .I1(n12320), .I2(n9759), .O(n7695) );
  ND2DHD U8806 ( .I1(n13821), .I2(n12089), .O(n11722) );
  ND3CHD U8807 ( .I1(n11874), .I2(n11873), .I3(n6851), .O(n10108) );
  ND2HHD U8808 ( .I1(n11873), .I2(n7389), .O(n11871) );
  NR2EHD U8809 ( .I1(n8371), .I2(n7879), .O(n10124) );
  ND2KHD U8810 ( .I1(n13653), .I2(n8628), .O(n8533) );
  INVQHD U8811 ( .I(n7841), .O(n7292) );
  AN2KHD U8812 ( .I1(n7788), .I2(n12086), .O(n12297) );
  ND2HHD U8813 ( .I1(n7859), .I2(n13659), .O(n8815) );
  ND3CHD U8814 ( .I1(n9612), .I2(n13821), .I3(n13659), .O(n11783) );
  ND3CHD U8815 ( .I1(n9612), .I2(n12302), .I3(n13659), .O(n9926) );
  NR2GHD U8816 ( .I1(n7148), .I2(n11838), .O(n11856) );
  OR3EHD U8817 ( .I1(n14086), .I2(n14085), .I3(n14084), .O(n14088) );
  NR2EHD U8818 ( .I1(n13243), .I2(n14084), .O(n8147) );
  NR2EHD U8819 ( .I1(n9357), .I2(n14084), .O(n9356) );
  OR2HHD U8820 ( .I1(n8754), .I2(n8753), .O(n7689) );
  ND2HHD U8821 ( .I1(n7219), .I2(_i_CLEFIA128_keyK _50), .O(n11672) );
  OA12HHD U8822 ( .B1(n9069), .B2(n8054), .A1(n14076), .O(n8053) );
  ND2KHD U8823 ( .I1(n9129), .I2(n10583), .O(n10568) );
  INVKHD U8824 ( .I(n10568), .O(n7081) );
  ND2HHD U8825 ( .I1(n7153), .I2(n10163), .O(n10162) );
  NR2GHD U8826 ( .I1(n13549), .I2(n11792), .O(n11800) );
  ND2KHD U8827 ( .I1(n11713), .I2(n7035), .O(n13506) );
  INVMHD U8828 ( .I(n13593), .O(n8184) );
  NR2IHD U8829 ( .I1(n7540), .I2(n8665), .O(n8717) );
  XNR2KHD U8830 ( .I1(n10460), .I2(n8741), .O(n6832) );
  XNR2KHD U8831 ( .I1(n10460), .I2(n8741), .O(n6833) );
  ND2KHD U8832 ( .I1(n6869), .I2(n9790), .O(n8741) );
  BUFKHD U8833 ( .I(n7998), .O(n7970) );
  NR2EHD U8834 ( .I1(n10860), .I2(n6906), .O(n10868) );
  ND3EHD U8835 ( .I1(n12735), .I2(n12725), .I3(n8462), .O(n8461) );
  NR2CHD U8836 ( .I1(n12671), .I2(n8563), .O(n8562) );
  INVKHD U8837 ( .I(n12793), .O(n8563) );
  INVNHD U8838 ( .I(n9366), .O(n9613) );
  ND2DHD U8839 ( .I1(n7316), .I2(n9007), .O(n9691) );
  ND3EHD U8840 ( .I1(n6918), .I2(n13629), .I3(n13125), .O(n13127) );
  NR2IHD U8841 ( .I1(n10633), .I2(n10634), .O(n7508) );
  ND2HHD U8842 ( .I1(n7185), .I2(n12651), .O(n10633) );
  ND2HHD U8843 ( .I1(n10269), .I2(n12646), .O(n7197) );
  ND2KHD U8844 ( .I1(n8226), .I2(n11818), .O(n14051) );
  ND2HHD U8845 ( .I1(n9538), .I2(n14696), .O(n14704) );
  NR2CHD U8846 ( .I1(n7959), .I2(n12271), .O(n7958) );
  OR2B1HHD U8847 ( .I1(n13576), .B1(n13122), .O(n12936) );
  AN3HHD U8848 ( .I1(n10823), .I2(n12687), .I3(n10822), .O(n9851) );
  INVMHD U8849 ( .I(n12864), .O(n12717) );
  OAI112EHD U8850 ( .C1(n13277), .C2(n15404), .A1(n13355), .B1(n13354), .O(n6307) );
  ND2DHD U8851 ( .I1(n15067), .I2(n11130), .O(n9616) );
  XNR2KHD U8852 ( .I1(_i_CLEFIA128_CON_T_x _1), .I2(DOUT_97), .O(n6834) );
  INVCKLHD U8853 ( .I(n8986), .O(n10169) );
  ND3HHD U8854 ( .I1(n12618), .I2(n12619), .I3(n12617), .O(n12625) );
  INVCKLHD U8855 ( .I(n10657), .O(n7347) );
  NR2CHD U8856 ( .I1(n8488), .I2(n11218), .O(n8487) );
  NR2CHD U8857 ( .I1(n12626), .I2(n10866), .O(n10867) );
  NR2GHD U8858 ( .I1(n11059), .I2(n11058), .O(n11201) );
  NR2EHD U8859 ( .I1(n12625), .I2(n10264), .O(n12631) );
  INVQHD U8860 ( .I(n6836), .O(n6837) );
  ND2HHD U8861 ( .I1(n9557), .I2(n9858), .O(n6838) );
  ND2HHD U8862 ( .I1(n9557), .I2(n9858), .O(n9912) );
  ND2HHD U8863 ( .I1(n9704), .I2(n12605), .O(n10270) );
  MUX2HHD U8864 ( .A(n10346), .B(n10345), .S(_i_CLEFIA128_keyL _95), .O(n10351) );
  ND3EHD U8865 ( .I1(n7187), .I2(n11079), .I3(n11250), .O(n12626) );
  NR3HHD U8866 ( .I1(n13490), .I2(n12186), .I3(n12183), .O(n9358) );
  ND2HHD U8867 ( .I1(n7187), .I2(n7359), .O(n11080) );
  NR2IHD U8868 ( .I1(n9566), .I2(n9565), .O(n8800) );
  INVJHD U8869 ( .I(n9191), .O(n10836) );
  ND2KHD U8870 ( .I1(n9676), .I2(n9430), .O(n13036) );
  XNR2KHD U8871 ( .I1(n14636), .I2(n13743), .O(n15152) );
  OAI12EHD U8872 ( .B1(n13432), .B2(n9214), .A1(n13440), .O(n9212) );
  ND2HHD U8873 ( .I1(n9595), .I2(n8451), .O(n9617) );
  NR2EHD U8874 ( .I1(n8118), .I2(n7484), .O(n9754) );
  INVGHD U8875 ( .I(n6844), .O(n6845) );
  ND2KHD U8876 ( .I1(n6819), .I2(n12766), .O(n11475) );
  XNR2HHD U8877 ( .I1(n10196), .I2(n10195), .O(n14938) );
  ND2HHD U8878 ( .I1(n8943), .I2(n7521), .O(n7520) );
  ND3EHD U8879 ( .I1(n14178), .I2(n14179), .I3(n14177), .O(n6179) );
  ND2DHD U8880 ( .I1(n9817), .I2(n11130), .O(n14178) );
  OR3HHD U8881 ( .I1(n10674), .I2(n10675), .I3(n10676), .O(n10677) );
  AN2EHD U8882 ( .I1(n11818), .I2(n6801), .O(n7702) );
  ND2HHD U8883 ( .I1(n12127), .I2(n12121), .O(n13143) );
  ND2HHD U8884 ( .I1(n8208), .I2(n6803), .O(n10844) );
  INVNHD U8885 ( .I(n12768), .O(n12752) );
  AN3HHD U8886 ( .I1(n12754), .I2(n12753), .I3(n12752), .O(n12755) );
  ND3EHD U8887 ( .I1(n12743), .I2(n12768), .I3(n12742), .O(n12745) );
  ND2DHD U8888 ( .I1(n12622), .I2(n12623), .O(n10265) );
  ND2HHD U8889 ( .I1(n10307), .I2(n6851), .O(n10309) );
  NR2EHD U8890 ( .I1(n11928), .I2(n9929), .O(n12991) );
  ND2KHD U8891 ( .I1(n7979), .I2(n7978), .O(n7972) );
  ND2KHD U8892 ( .I1(n7320), .I2(n7319), .O(n7302) );
  AN3EHD U8893 ( .I1(n12610), .I2(n6803), .I3(n11250), .O(n11251) );
  AN2EHD U8894 ( .I1(n9460), .I2(n6803), .O(n10770) );
  BUFQHD U8895 ( .I(n11999), .O(n12915) );
  XNR2KHD U8896 ( .I1(_i_CLEFIA128_CON_T_x _14), .I2(DOUT_61), .O(n8447) );
  ND2HHD U8897 ( .I1(n10465), .I2(n6851), .O(n10242) );
  BUFQHD U8898 ( .I(n12118), .O(n10095) );
  BUFQHD U8899 ( .I(n7574), .O(n6843) );
  ND3CHD U8900 ( .I1(n12502), .I2(n6894), .I3(n11300), .O(n11302) );
  ND2HHD U8901 ( .I1(n11865), .I2(n6845), .O(n11867) );
  INVQHD U8902 ( .I(_i_CLEFIA128_keyL _40), .O(n15281) );
  ND2HHD U8903 ( .I1(n9175), .I2(n6851), .O(n9171) );
  NR2IHD U8904 ( .I1(n8798), .I2(n8173), .O(n8174) );
  INVQHD U8905 ( .I(_i_CLEFIA128_keyK _93), .O(n8173) );
  NR2EHD U8906 ( .I1(n7626), .I2(n7623), .O(n7622) );
  NR2EHD U8907 ( .I1(n11111), .I2(n8473), .O(n8472) );
  ND2KHD U8908 ( .I1(n11948), .I2(n7830), .O(n13425) );
  AN2KHD U8909 ( .I1(n13425), .I2(n10295), .O(n9216) );
  ND2KHD U8910 ( .I1(n11930), .I2(n11904), .O(n11893) );
  ND3EHD U8911 ( .I1(n10212), .I2(n13242), .I3(n13241), .O(n7921) );
  BUFMHD U8912 ( .I(n11245), .O(n6846) );
  ND2HHD U8913 ( .I1(n9950), .I2(n6851), .O(n7328) );
  NR2EHD U8914 ( .I1(n7167), .I2(n8456), .O(n8455) );
  BUFMHD U8915 ( .I(n8452), .O(n8018) );
  NR2GHD U8916 ( .I1(n11572), .I2(n14707), .O(n10190) );
  ND2HHD U8917 ( .I1(n14083), .I2(n14056), .O(n13253) );
  NR2IHD U8918 ( .I1(n11647), .I2(n11832), .O(n14059) );
  ND2DHD U8919 ( .I1(n6682), .I2(n13643), .O(n13644) );
  ND2HHD U8920 ( .I1(n8723), .I2(n8563), .O(n8722) );
  OAI13HHD U8921 ( .B1(n12787), .B2(n12786), .B3(n12785), .A1(n10282), .O(n8985) );
  INVKHD U8922 ( .I(n12685), .O(n10282) );
  ND2DHD U8923 ( .I1(n7104), .I2(n10687), .O(n6847) );
  ND2HHD U8924 ( .I1(n12764), .I2(n6849), .O(n9610) );
  ND3EHD U8925 ( .I1(n12640), .I2(n8235), .I3(n8208), .O(n7127) );
  ND3EHD U8926 ( .I1(n8264), .I2(n13444), .I3(n13443), .O(n13445) );
  NR2EHD U8927 ( .I1(n13446), .I2(n13445), .O(n13452) );
  ND3EHD U8928 ( .I1(n13453), .I2(n13452), .I3(n13451), .O(n13455) );
  INVQHD U8929 ( .I(n6850), .O(n6851) );
  INVKHD U8930 ( .I(n7138), .O(n8220) );
  ND3CHD U8931 ( .I1(n9909), .I2(n12357), .I3(n7561), .O(n9889) );
  NR2IHD U8932 ( .I1(n8128), .I2(n8129), .O(n8127) );
  AN2KHD U8933 ( .I1(n13241), .I2(n13216), .O(n14067) );
  AN2EHD U8934 ( .I1(n10193), .I2(n14076), .O(n8414) );
  ND2DHD U8935 ( .I1(n9564), .I2(n14076), .O(n9227) );
  OA12EHD U8936 ( .B1(n14077), .B2(n7713), .A1(n14076), .O(n7712) );
  INVGHD U8937 ( .I(n7414), .O(n7412) );
  ND2HHD U8938 ( .I1(n10680), .I2(n12603), .O(n10682) );
  ND2DHD U8939 ( .I1(_i_CLEFIA128_keyL _49), .I2(n7219), .O(n8660) );
  INVGHD U8940 ( .I(n8763), .O(n8166) );
  ND2HHD U8941 ( .I1(n8763), .I2(n10107), .O(n8114) );
  ND3EHD U8942 ( .I1(n11862), .I2(n14405), .I3(_i_CLEFIA128_keyL _108), .O(n11863) );
  OR2KHD U8943 ( .I1(n11612), .I2(n9493), .O(n8760) );
  NR2IHD U8944 ( .I1(n9481), .I2(n9480), .O(n9479) );
  ND3EHD U8945 ( .I1(n10051), .I2(n6931), .I3(n6831), .O(n9481) );
  INVQHD U8946 ( .I(_i_CLEFIA128_keyL _99), .O(n15404) );
  INVNHD U8947 ( .I(n12497), .O(n10720) );
  ND2DHD U8948 ( .I1(n9567), .I2(n8995), .O(n6852) );
  NR2IHD U8949 ( .I1(n12408), .I2(n12409), .O(n8995) );
  NR2IHD U8950 ( .I1(n9602), .I2(n9860), .O(n9567) );
  OA112HHD U8951 ( .C1(n11275), .C2(n11285), .A1(n9012), .B1(n12450), .O(n11278) );
  INVQHD U8952 ( .I(n9541), .O(n9626) );
  INVNHD U8953 ( .I(n8739), .O(n9541) );
  NR2IHD U8954 ( .I1(n11559), .I2(n11539), .O(n9105) );
  ND2HHD U8955 ( .I1(n6873), .I2(n12484), .O(n9135) );
  ND3EHD U8956 ( .I1(n6853), .I2(n6855), .I3(n6854), .O(n6856) );
  AN2HHD U8957 ( .I1(n6856), .I2(n12462), .O(n9052) );
  ND3EHD U8958 ( .I1(n11314), .I2(n11278), .I3(n11277), .O(n11281) );
  XNR2KHD U8959 ( .I1(n14996), .I2(n10161), .O(n9930) );
  OR3HHD U8960 ( .I1(n12300), .I2(n11726), .I3(n11803), .O(n11728) );
  NR2IHD U8961 ( .I1(n7236), .I2(n7235), .O(n9643) );
  OA13EHD U8962 ( .B1(n11527), .B2(n11536), .B3(n11528), .A1(n12474), .O(n11540) );
  BUFQHD U8963 ( .I(n8589), .O(n7389) );
  OR3EHD U8964 ( .I1(n9436), .I2(n13362), .I3(n9672), .O(n13363) );
  NR2IHD U8965 ( .I1(n8179), .I2(n7209), .O(n10570) );
  INVQHD U8966 ( .I(n6884), .O(n11911) );
  ND2DHD U8967 ( .I1(n13036), .I2(n9093), .O(n12229) );
  AN2EHD U8968 ( .I1(n13401), .I2(n13036), .O(n12951) );
  ND2DHD U8969 ( .I1(n10459), .I2(n8589), .O(n7649) );
  ND2KHD U8970 ( .I1(n12497), .I2(n10617), .O(n9256) );
  XOR2EHD U8971 ( .I1(n14328), .I2(n14329), .O(n14634) );
  ND2DHD U8972 ( .I1(n7002), .I2(n11446), .O(n11451) );
  AN2EHD U8973 ( .I1(n7376), .I2(n11295), .O(n7378) );
  NR2GHD U8974 ( .I1(n7040), .I2(n7209), .O(n11416) );
  NR2GHD U8975 ( .I1(n9100), .I2(n6859), .O(n6858) );
  ND2DHD U8976 ( .I1(n11429), .I2(n12478), .O(n6859) );
  INVHHD U8977 ( .I(n9100), .O(n9238) );
  ND2HHD U8978 ( .I1(n11297), .I2(n12453), .O(n9100) );
  INVNHD U8979 ( .I(n8850), .O(n11906) );
  ND2HHD U8980 ( .I1(n6863), .I2(n6862), .O(n6861) );
  AN2HHD U8981 ( .I1(n9842), .I2(n11503), .O(n6862) );
  ND3CHD U8982 ( .I1(n13251), .I2(n7967), .I3(n7842), .O(n13252) );
  AN2EHD U8983 ( .I1(n7842), .I2(n13085), .O(n11641) );
  BUFQHD U8984 ( .I(n11631), .O(n8210) );
  NR2IHD U8985 ( .I1(n11540), .I2(n11560), .O(n9066) );
  ND2KHD U8986 ( .I1(n8343), .I2(n12476), .O(n6865) );
  ND2KHD U8987 ( .I1(n9288), .I2(n6866), .O(n9287) );
  INVKHD U8988 ( .I(n6865), .O(n6866) );
  ND3CHD U8989 ( .I1(n12094), .I2(n13673), .I3(n9405), .O(n12095) );
  ND3CHD U8990 ( .I1(n13396), .I2(n13371), .I3(n9847), .O(n9911) );
  ND2HHD U8991 ( .I1(n11498), .I2(n11499), .O(n11501) );
  ND2KHD U8992 ( .I1(n12056), .I2(n9580), .O(n8729) );
  ND2DHD U8993 ( .I1(n7398), .I2(n9694), .O(n6867) );
  ND3CHD U8994 ( .I1(n11840), .I2(n9184), .I3(n9568), .O(n11841) );
  INVNHD U8995 ( .I(n10208), .O(n12216) );
  NR2GHD U8996 ( .I1(n12962), .I2(n9620), .O(n9642) );
  ND3CHD U8997 ( .I1(n11845), .I2(n13483), .I3(n7594), .O(n11846) );
  NR2EHD U8998 ( .I1(n12757), .I2(n10529), .O(n10531) );
  INVNHD U8999 ( .I(n8780), .O(n12424) );
  ND2HHD U9000 ( .I1(n7383), .I2(n6931), .O(n11811) );
  NR2IHD U9001 ( .I1(n7808), .I2(n8083), .O(n11794) );
  ND3EHD U9002 ( .I1(n7118), .I2(n8197), .I3(n13083), .O(n13054) );
  ND2HHD U9003 ( .I1(n11628), .I2(n11612), .O(n11762) );
  AN2EHD U9004 ( .I1(n12124), .I2(n8729), .O(n10186) );
  BUFMHD U9005 ( .I(n11677), .O(n13521) );
  ND2DHD U9006 ( .I1(n14913), .I2(n11130), .O(n13564) );
  OR2HHD U9007 ( .I1(n9525), .I2(n12168), .O(n7121) );
  INVDHD U9008 ( .I(n9799), .O(n9360) );
  BUFEHD U9009 ( .I(n7943), .O(n7935) );
  ND2HHD U9010 ( .I1(n6694), .I2(n7859), .O(n11782) );
  NR2EHD U9011 ( .I1(n11804), .I2(n9001), .O(n8652) );
  INVMHD U9012 ( .I(n11904), .O(n7811) );
  XNR2KHD U9013 ( .I1(n14109), .I2(n9370), .O(n14184) );
  NR2GHD U9014 ( .I1(n9156), .I2(n9371), .O(n14109) );
  INVNHD U9015 ( .I(n10252), .O(n6873) );
  ND2HHD U9016 ( .I1(n14342), .I2(n14343), .O(n9371) );
  ND2DHD U9017 ( .I1(n14343), .I2(n14342), .O(n7927) );
  ND2HHD U9018 ( .I1(n7928), .I2(n13826), .O(n14342) );
  ND2HHD U9019 ( .I1(n14913), .I2(n14886), .O(n14894) );
  XNR2EHD U9020 ( .I1(n14109), .I2(n9776), .O(n14031) );
  ND2HHD U9021 ( .I1(n12163), .I2(n12162), .O(n13645) );
  NR2GHD U9022 ( .I1(n13645), .I2(n12164), .O(n12165) );
  ND2HHD U9023 ( .I1(n12304), .I2(n8538), .O(n7427) );
  NR2GHD U9024 ( .I1(n8539), .I2(n8540), .O(n8538) );
  NR2IHD U9025 ( .I1(n7700), .I2(n11778), .O(n11781) );
  ND3CHD U9026 ( .I1(n7619), .I2(n8589), .I3(_i_CLEFIA128_keyL _82), .O(n7618) );
  XOR2CHD U9027 ( .I1(n7557), .I2(_i_CLEFIA128_keyL _96), .O(n6886) );
  XOR2EHD U9028 ( .I1(n6852), .I2(n14108), .O(n10127) );
  NR2GHD U9029 ( .I1(n10021), .I2(n7826), .O(n7829) );
  ND2HHD U9030 ( .I1(n11648), .I2(n7044), .O(n6875) );
  XNR2KHD U9031 ( .I1(n6877), .I2(n7549), .O(n7547) );
  NR2EHD U9032 ( .I1(n7949), .I2(n8890), .O(n7948) );
  NR2IHD U9033 ( .I1(n7653), .I2(n7651), .O(n7087) );
  XNR2HHD U9034 ( .I1(n15120), .I2(n11983), .O(n6878) );
  XNR2HHD U9035 ( .I1(n15120), .I2(n11983), .O(n11985) );
  ND2DHD U9036 ( .I1(n9992), .I2(n10959), .O(n8145) );
  AN2HHD U9037 ( .I1(n12302), .I2(n8581), .O(n10036) );
  INVGHD U9038 ( .I(n9415), .O(n6880) );
  ND2HHD U9039 ( .I1(n8101), .I2(n10485), .O(n8100) );
  AN3EHD U9040 ( .I1(n11512), .I2(n10485), .I3(n11511), .O(n11513) );
  BUFQHD U9041 ( .I(n12066), .O(n9807) );
  INVMHD U9042 ( .I(n9701), .O(n11996) );
  ND2KHD U9043 ( .I1(n9742), .I2(n9667), .O(n11616) );
  ND2HHD U9044 ( .I1(n8865), .I2(n8864), .O(n14138) );
  AN2HHD U9045 ( .I1(n11411), .I2(n6621), .O(n8387) );
  NR2IHD U9046 ( .I1(n10669), .I2(n9261), .O(n8983) );
  AN2EHD U9047 ( .I1(n12163), .I2(n12302), .O(n8299) );
  ND3CHD U9048 ( .I1(n12655), .I2(n9145), .I3(n11079), .O(n7322) );
  ND3EHD U9049 ( .I1(n8039), .I2(n9528), .I3(_i_CLEFIA128_keyK _73), .O(n8945) );
  ND2KHD U9050 ( .I1(n13471), .I2(n7967), .O(n9695) );
  ND2DHD U9051 ( .I1(n14433), .I2(_i_CLEFIA128_CON_T_x _1), .O(n14750) );
  INVCKGHD U9052 ( .I(n10085), .O(n9902) );
  AN2HHD U9053 ( .I1(n8115), .I2(n10051), .O(n6938) );
  NR2EHD U9054 ( .I1(n10902), .I2(n10901), .O(n10903) );
  INVMHD U9055 ( .I(n7977), .O(n11840) );
  BUFQHD U9056 ( .I(n10293), .O(n9581) );
  ND2KHD U9057 ( .I1(n8196), .I2(n7810), .O(n8583) );
  NR2IHD U9058 ( .I1(n10051), .I2(n8083), .O(n8992) );
  NR2EHD U9059 ( .I1(n12670), .I2(n8968), .O(n8967) );
  ND2KHD U9060 ( .I1(n8200), .I2(n7933), .O(n13646) );
  NR2CHD U9061 ( .I1(n13243), .I2(n11767), .O(n11768) );
  XNR2KHD U9062 ( .I1(n6885), .I2(n8675), .O(n6884) );
  INVNHD U9063 ( .I(n8115), .O(n9830) );
  ND2DHD U9064 ( .I1(n9455), .I2(n7336), .O(n14044) );
  AO12HHD U9065 ( .B1(n10154), .B2(n13112), .A1(n9536), .O(n10153) );
  ND3HHD U9066 ( .I1(n7165), .I2(n9832), .I3(n13595), .O(n13192) );
  ND2DHD U9067 ( .I1(n12604), .I2(n12603), .O(n12606) );
  ND3CHD U9068 ( .I1(n10366), .I2(n12603), .I3(n8911), .O(n10367) );
  INVGHD U9069 ( .I(n13642), .O(n9155) );
  ND2DHD U9070 ( .I1(n12299), .I2(n13642), .O(n11725) );
  INVJHD U9071 ( .I(n13014), .O(n9081) );
  ND3HHD U9072 ( .I1(n9621), .I2(n12150), .I3(n12065), .O(n12068) );
  ND2KHD U9073 ( .I1(n7772), .I2(n8952), .O(n7234) );
  ND2HHD U9074 ( .I1(n15024), .I2(n15002), .O(n15010) );
  AN3HHD U9075 ( .I1(n12688), .I2(n12690), .I3(n8914), .O(n6915) );
  XNR2KHD U9076 ( .I1(n8068), .I2(n8067), .O(n6887) );
  INVQHD U9077 ( .I(_i_CLEFIA128_keyL _80), .O(n8902) );
  ND3EHD U9078 ( .I1(n6997), .I2(n9708), .I3(n10022), .O(n6888) );
  NR2EHD U9079 ( .I1(n7466), .I2(n7465), .O(n7464) );
  ND2HHD U9080 ( .I1(n9882), .I2(n13608), .O(n9881) );
  ND2DHD U9081 ( .I1(n11175), .I2(n11176), .O(n12487) );
  NR2CHD U9082 ( .I1(n11279), .I2(n10975), .O(n10983) );
  INVGHD U9083 ( .I(n8930), .O(n8929) );
  NR2EHD U9084 ( .I1(n8930), .I2(n8616), .O(n10416) );
  ND2HHD U9085 ( .I1(n6716), .I2(n8495), .O(n12780) );
  INVJHD U9086 ( .I(n12592), .O(n7021) );
  ND2KHD U9087 ( .I1(n9694), .I2(n8182), .O(n11382) );
  XOR2HHD U9088 ( .I1(_i_CLEFIA128_CON_T_x _6), .I2(DOUT_45), .O(n10417) );
  XNR2KHD U9089 ( .I1(n6890), .I2(n8717), .O(n11680) );
  ND2DHD U9090 ( .I1(n8657), .I2(n12268), .O(n7463) );
  ND3HHD U9091 ( .I1(n13614), .I2(n13613), .I3(n13612), .O(n13616) );
  XOR2HHD U9092 ( .I1(_i_CLEFIA128_keyL _100), .I2(n11964), .O(n11965) );
  AN2HHD U9093 ( .I1(n12553), .I2(n7539), .O(n6947) );
  XNR2KHD U9094 ( .I1(n14230), .I2(n14229), .O(n15054) );
  NR2EHD U9095 ( .I1(n8897), .I2(n6810), .O(n12901) );
  BUFNHD U9096 ( .I(n9635), .O(n8881) );
  NR2EHD U9097 ( .I1(n11451), .I2(n11450), .O(n11456) );
  NR2EHD U9098 ( .I1(n12573), .I2(n12576), .O(n7277) );
  INVNHD U9099 ( .I(n10325), .O(n10659) );
  ND2HHD U9100 ( .I1(n8521), .I2(n15500), .O(n9788) );
  INVNHD U9101 ( .I(n8778), .O(n9684) );
  INVMHD U9102 ( .I(n11685), .O(n10266) );
  ND2KHD U9103 ( .I1(n13659), .I2(n12299), .O(n8856) );
  NR2CHD U9104 ( .I1(n12294), .I2(n9070), .O(n7511) );
  INVCKGHD U9105 ( .I(n13183), .O(n10128) );
  ND2KHD U9106 ( .I1(n9772), .I2(n8866), .O(n7409) );
  XNR2KHD U9107 ( .I1(n6924), .I2(n7390), .O(n12349) );
  ND2KHD U9108 ( .I1(n7598), .I2(n7601), .O(n13972) );
  NR2IHD U9109 ( .I1(n7600), .I2(n7599), .O(n7598) );
  ND2KHD U9110 ( .I1(n9903), .I2(n9800), .O(n12469) );
  INVNHD U9111 ( .I(n12500), .O(n6892) );
  INVNHD U9112 ( .I(n6892), .O(n6894) );
  ND2DHD U9113 ( .I1(n8235), .I2(n12537), .O(n10386) );
  INVJHD U9114 ( .I(n8182), .O(n11324) );
  INVQHD U9115 ( .I(n8181), .O(n8182) );
  NR2IHD U9116 ( .I1(n7799), .I2(n7798), .O(n9547) );
  ND2KHD U9117 ( .I1(n11943), .I2(n11948), .O(n7393) );
  XNR2KHD U9118 ( .I1(_i_CLEFIA128_keyL _114), .I2(n8122), .O(n11675) );
  NR2GHD U9119 ( .I1(n8477), .I2(n12759), .O(n8475) );
  NR2EHD U9120 ( .I1(n13816), .I2(n13808), .O(n7845) );
  INVGHD U9121 ( .I(n12297), .O(n7670) );
  ND2HHD U9122 ( .I1(n12297), .I2(n13684), .O(n7615) );
  ND2DHD U9123 ( .I1(n12066), .I2(n7773), .O(n11813) );
  ND2HHD U9124 ( .I1(n9040), .I2(n13622), .O(n9880) );
  ND2DHD U9125 ( .I1(n11403), .I2(n11360), .O(n11321) );
  INVNHD U9126 ( .I(n7756), .O(n8215) );
  ND2HHD U9127 ( .I1(n8039), .I2(_i_CLEFIA128_keyK _10), .O(n10407) );
  INVCKIHD U9128 ( .I(n7451), .O(n7521) );
  BUFQHD U9129 ( .I(n11794), .O(n7809) );
  BUFHHD U9130 ( .I(n12520), .O(n7128) );
  NR2EHD U9131 ( .I1(n10377), .I2(n11264), .O(n10378) );
  ND2HHD U9132 ( .I1(n10849), .I2(n12652), .O(n11264) );
  INVNHD U9133 ( .I(n10481), .O(n9841) );
  INVLHD U9134 ( .I(n12512), .O(n7344) );
  ND2HHD U9135 ( .I1(_i_CLEFIA128_keyK _1), .I2(_i_CLEFIA128_keyL _1), .O(n10463) );
  NR2CHD U9136 ( .I1(n7377), .I2(n11165), .O(n11174) );
  ND3CHD U9137 ( .I1(n11256), .I2(n11255), .I3(n7178), .O(n11257) );
  NR2EHD U9138 ( .I1(n11257), .I2(n11258), .O(n11267) );
  INVJHD U9139 ( .I(n6864), .O(n7673) );
  ND2HHD U9140 ( .I1(n13821), .I2(n13842), .O(n11714) );
  NR2IHD U9141 ( .I1(n12400), .I2(n12399), .O(n13120) );
  OAI22EHD U9142 ( .A1(n12561), .A2(n8116), .B1(n9050), .B2(n8182), .O(n12563));
  AN2HHD U9143 ( .I1(n12501), .I2(n11541), .O(n11188) );
  OR3EHD U9144 ( .I1(n9728), .I2(n12058), .I3(n7488), .O(n9979) );
  NR2IHD U9145 ( .I1(n12260), .I2(n12261), .O(n12274) );
  NR2IHD U9146 ( .I1(n9036), .I2(n11471), .O(n10043) );
  AN2EHD U9147 ( .I1(n10251), .I2(n12501), .O(n8769) );
  ND3CHD U9148 ( .I1(n11522), .I2(n11429), .I3(n12501), .O(n11453) );
  ND2HHD U9149 ( .I1(n8767), .I2(n10973), .O(n11443) );
  OAI12EHD U9150 ( .B1(n15054), .B2(n15416), .A1(n14585), .O(n6284) );
  INVJHD U9151 ( .I(n12226), .O(n11908) );
  ND2HHD U9152 ( .I1(n7900), .I2(n12448), .O(n12494) );
  XOR2EHD U9153 ( .I1(n14352), .I2(n14228), .O(n14229) );
  ND2DHD U9154 ( .I1(n9721), .I2(n9175), .O(n9172) );
  INVGHD U9155 ( .I(n7673), .O(n6896) );
  ND2DHD U9156 ( .I1(n7597), .I2(n10760), .O(n9523) );
  NR2GHD U9157 ( .I1(n10472), .I2(n9750), .O(n10473) );
  ND2DHD U9158 ( .I1(n12502), .I2(n6894), .O(n7273) );
  NR2IHD U9159 ( .I1(n13669), .I2(n13668), .O(n9820) );
  NR2GHD U9160 ( .I1(n11085), .I2(n7344), .O(n7323) );
  ND2KHD U9161 ( .I1(n13194), .I2(n13629), .O(n10129) );
  BUFQHD U9162 ( .I(n8227), .O(n7907) );
  NR2EHD U9163 ( .I1(n13068), .I2(n13067), .O(n13070) );
  INVGHD U9164 ( .I(n12123), .O(n13172) );
  ND2HHD U9165 ( .I1(n13121), .I2(n12123), .O(n7469) );
  ND3CHD U9166 ( .I1(n13128), .I2(n12123), .I3(n13572), .O(n10013) );
  ND2KHD U9167 ( .I1(n9855), .I2(n7597), .O(n12847) );
  ND3CHD U9168 ( .I1(n11015), .I2(n11014), .I3(n11360), .O(n11016) );
  ND2KHD U9169 ( .I1(n8191), .I2(n8215), .O(n8979) );
  OA12EHD U9170 ( .B1(n15404), .B2(_i_CLEFIA128_keyK _99), .A1(n14405), .O(n11968) );
  ND2DHD U9171 ( .I1(n10550), .I2(n6851), .O(n7914) );
  ND2DHD U9172 ( .I1(n10030), .I2(n6851), .O(n10029) );
  NR2IHD U9173 ( .I1(n9975), .I2(n7733), .O(n12854) );
  INVNHD U9174 ( .I(n12029), .O(n10228) );
  ND2HHD U9175 ( .I1(n12902), .I2(n10095), .O(n13603) );
  ND2KHD U9176 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(n8797), .O(n6898) );
  ND2KHD U9177 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(n8797), .O(n6899) );
  ND3EHD U9178 ( .I1(n8987), .I2(n7878), .I3(n7877), .O(n6900) );
  BUFKHD U9179 ( .I(n14707), .O(n7103) );
  ND2KHD U9180 ( .I1(n13053), .I2(n8026), .O(n12196) );
  INVJHD U9181 ( .I(n10326), .O(n10636) );
  INVJHD U9182 ( .I(n6902), .O(n6903) );
  NR2EHD U9183 ( .I1(n8458), .I2(n8461), .O(n8457) );
  INVJHD U9184 ( .I(n12585), .O(n9352) );
  INVCKGHD U9185 ( .I(n8595), .O(n7421) );
  ND2HHD U9186 ( .I1(n9356), .I2(n9358), .O(n9445) );
  NR2GHD U9187 ( .I1(n10385), .I2(n10386), .O(n10859) );
  ND2DHD U9188 ( .I1(n7359), .I2(n9344), .O(n10385) );
  NR2EHD U9189 ( .I1(n12196), .I2(n13489), .O(n8025) );
  INVQHD U9190 ( .I(n8219), .O(n9811) );
  INVNHD U9191 ( .I(n7105), .O(n8219) );
  INVMHD U9192 ( .I(n7458), .O(n8115) );
  XNR3EHD U9193 ( .I1(n10262), .I2(n14636), .I3(n9743), .O(n6904) );
  XOR2KHD U9194 ( .I1(n9923), .I2(n10149), .O(n14636) );
  ND2DHD U9195 ( .I1(n12190), .I2(n11763), .O(n9510) );
  ND2DHD U9196 ( .I1(n7704), .I2(n9186), .O(n12191) );
  AN2EHD U9197 ( .I1(n11911), .I2(n7811), .O(n6930) );
  ND2HHD U9198 ( .I1(n12677), .I2(n10964), .O(n10285) );
  NR2GHD U9199 ( .I1(n7526), .I2(n7525), .O(n7524) );
  INVMHD U9200 ( .I(n7776), .O(n7198) );
  BUFQHD U9201 ( .I(n7930), .O(n7254) );
  ND2KHD U9202 ( .I1(n9807), .I2(n7254), .O(n9152) );
  ND2HHD U9203 ( .I1(n9531), .I2(n11552), .O(n8094) );
  ND3EHD U9204 ( .I1(n13071), .I2(n13069), .I3(n13070), .O(n13074) );
  NR2EHD U9205 ( .I1(n8998), .I2(n8997), .O(n8996) );
  ND2DHD U9206 ( .I1(n12179), .I2(n10146), .O(n8762) );
  INVJHD U9207 ( .I(n9661), .O(n12676) );
  ND2HHD U9208 ( .I1(n8977), .I2(n10945), .O(n9661) );
  ND2HHD U9209 ( .I1(n8331), .I2(n13478), .O(n8084) );
  INVJHD U9210 ( .I(n7700), .O(n13833) );
  ND2DHD U9211 ( .I1(n7779), .I2(n12522), .O(n11064) );
  ND2DHD U9212 ( .I1(n8208), .I2(n7779), .O(n12539) );
  XNR2KHD U9213 ( .I1(n9442), .I2(n7479), .O(n6905) );
  ND3EHD U9214 ( .I1(n6992), .I2(n7122), .I3(n7183), .O(n6906) );
  INVQHD U9215 ( .I(n8798), .O(n7051) );
  INVQHD U9216 ( .I(n8798), .O(n8039) );
  ND2DHD U9217 ( .I1(n10990), .I2(n9627), .O(n11276) );
  ND2DHD U9218 ( .I1(n7671), .I2(n9626), .O(n8781) );
  ND2HHD U9219 ( .I1(n9626), .I2(n7671), .O(n9627) );
  XNR2HHD U9220 ( .I1(n6880), .I2(n14141), .O(n9938) );
  ND2HHD U9221 ( .I1(n9238), .I2(n11418), .O(n11422) );
  NR2IHD U9222 ( .I1(n7300), .I2(n7299), .O(n13107) );
  ND3EHD U9223 ( .I1(n11353), .I2(n12571), .I3(n11354), .O(n11355) );
  OA12HHD U9224 ( .B1(n12961), .B2(n12960), .A1(n13431), .O(n6907) );
  ND3EHD U9225 ( .I1(n12959), .I2(n9117), .I3(n12958), .O(n12960) );
  AN2HHD U9226 ( .I1(n8470), .I2(n11323), .O(n8469) );
  NR2EHD U9227 ( .I1(n13515), .I2(n13514), .O(n13516) );
  ND2KHD U9228 ( .I1(n11681), .I2(n12145), .O(n13651) );
  INVNHD U9229 ( .I(n7774), .O(n11681) );
  BUFQHD U9230 ( .I(n10420), .O(n10760) );
  NR2IHD U9231 ( .I1(n9859), .I2(n9861), .O(n9858) );
  INVNHD U9232 ( .I(n8165), .O(n8214) );
  NR2IHD U9233 ( .I1(n12196), .I2(n13243), .O(n7504) );
  NR2CHD U9234 ( .I1(n8207), .I2(n10441), .O(n10741) );
  XOR2HHD U9235 ( .I1(n6908), .I2(n13926), .O(n9915) );
  XNR2HHD U9236 ( .I1(DOUT_3), .I2(n7256), .O(n6908) );
  ND2HHD U9237 ( .I1(n12418), .I2(n12341), .O(n12342) );
  NR2EHD U9238 ( .I1(n12340), .I2(n12339), .O(n12341) );
  ND2HHD U9239 ( .I1(n10622), .I2(n10623), .O(n10694) );
  ND3CHD U9240 ( .I1(n7376), .I2(n9298), .I3(n9128), .O(n10620) );
  ND2HHD U9241 ( .I1(n10904), .I2(n8233), .O(n7448) );
  OR3HHD U9242 ( .I1(n11179), .I2(n11448), .I3(n10626), .O(n10627) );
  ND2DHD U9243 ( .I1(n10076), .I2(n7043), .O(n10044) );
  ND2DHD U9244 ( .I1(n10076), .I2(n11130), .O(n10204) );
  INVQHD U9245 ( .I(n8211), .O(n12498) );
  ND3CHD U9246 ( .I1(n12274), .I2(n12273), .I3(n7958), .O(n7957) );
  ND2HHD U9247 ( .I1(n7301), .I2(n9049), .O(n8454) );
  ND2DHD U9248 ( .I1(n12585), .I2(n12730), .O(n12588) );
  AN2HHD U9249 ( .I1(n13019), .I2(n12347), .O(n12968) );
  ND2HHD U9250 ( .I1(n14101), .I2(n14100), .O(n6134) );
  XNR3EHD U9251 ( .I1(n6910), .I2(n14245), .I3(n14244), .O(n7055) );
  XNR2EHD U9252 ( .I1(DOUT_5), .I2(n8756), .O(n6910) );
  NR2IHD U9253 ( .I1(n7294), .I2(n7293), .O(n12179) );
  OA13HHD U9254 ( .B1(n13825), .B2(n12167), .B3(n13663), .A1(n13817), .O(n7294) );
  NR2IHD U9255 ( .I1(n8319), .I2(n9169), .O(n7047) );
  XNR2HHD U9256 ( .I1(n10117), .I2(n10116), .O(n14837) );
  ND2KHD U9257 ( .I1(n10702), .I2(n10703), .O(n11467) );
  NR2GHD U9258 ( .I1(n11447), .I2(n10700), .O(n10703) );
  NR2IHD U9259 ( .I1(n11779), .I2(n8006), .O(n8611) );
  NR2GHD U9260 ( .I1(n7857), .I2(n10138), .O(n9414) );
  ND2DHD U9261 ( .I1(_i_CLEFIA128_keyK _12), .I2(_i_CLEFIA128_keyL _12), .O(n10410) );
  OA12EHD U9262 ( .B1(n8106), .B2(n8105), .A1(_i_CLEFIA128_state_reg _1), .O(n8104) );
  ND2DHD U9263 ( .I1(n8183), .I2(n12134), .O(n9888) );
  INVDHD U9264 ( .I(n11929), .O(n10106) );
  AN2EHD U9265 ( .I1(n9330), .I2(n6578), .O(n8225) );
  INVDHD U9266 ( .I(n12478), .O(n9138) );
  NR2EHD U9267 ( .I1(n11089), .I2(n9351), .O(n9350) );
  AN2EHD U9268 ( .I1(n10899), .I2(n8232), .O(n10900) );
  ND2HHD U9269 ( .I1(n7039), .I2(n8182), .O(n11496) );
  INVDHD U9270 ( .I(n12568), .O(n12560) );
  AN2EHD U9271 ( .I1(n13680), .I2(n13537), .O(n13539) );
  ND2DHD U9272 ( .I1(n9770), .I2(n8866), .O(n13117) );
  NR2GHD U9273 ( .I1(n11788), .I2(n8821), .O(n13526) );
  ND3CHD U9274 ( .I1(n6770), .I2(n12989), .I3(n12988), .O(n12990) );
  INVDHD U9275 ( .I(n12388), .O(n7555) );
  ND2HHD U9276 ( .I1(n11529), .I2(n9298), .O(n12457) );
  ND3CHD U9277 ( .I1(n12502), .I2(n12453), .I3(n6894), .O(n11273) );
  AN2EHD U9278 ( .I1(n7369), .I2(n9492), .O(n11835) );
  NR2CHD U9279 ( .I1(n8625), .I2(n10100), .O(n10099) );
  ND2DHD U9280 ( .I1(n13511), .I2(n8351), .O(n13518) );
  NR2EHD U9281 ( .I1(n11789), .I2(n11790), .O(n13530) );
  AN3B1EHD U9282 ( .I1(n9927), .I2(n8424), .B1(n8884), .O(n9248) );
  INVDHD U9283 ( .I(n13126), .O(n7556) );
  AN2EHD U9284 ( .I1(n12736), .I2(n11323), .O(n8338) );
  NR2CHD U9285 ( .I1(n10476), .I2(n9036), .O(n10477) );
  NR2CHD U9286 ( .I1(n10980), .I2(n10979), .O(n10981) );
  NR2EHD U9287 ( .I1(n12707), .I2(n12706), .O(n7823) );
  NR2EHD U9288 ( .I1(n11260), .I2(n11259), .O(n12615) );
  ND2DHD U9289 ( .I1(n8838), .I2(n8840), .O(n8837) );
  INVDHD U9290 ( .I(n9223), .O(n12489) );
  INVDHD U9291 ( .I(n11087), .O(n7519) );
  ND2DHD U9292 ( .I1(n12476), .I2(n10277), .O(n10276) );
  INVCKLHD U9293 ( .I(_i_CLEFIA128_keyK _107), .O(n11857) );
  INVKHD U9294 ( .I(_i_CLEFIA128_keyL _41), .O(n15124) );
  XOR2EHD U9295 ( .I1(DOUT_9), .I2(n8561), .O(n13754) );
  INVDHD U9296 ( .I(_i_CLEFIA128_keyL _39), .O(n9478) );
  INVKHD U9297 ( .I(_i_CLEFIA128_keyL _49), .O(n15150) );
  INVJHD U9298 ( .I(_i_CLEFIA128_keyL _4), .O(n14934) );
  INVDHD U9299 ( .I(_i_CLEFIA128_keyL _0), .O(n15146) );
  ND2DHD U9300 ( .I1(n7725), .I2(n11130), .O(n14175) );
  AN2HHD U9301 ( .I1(n12389), .I2(n7555), .O(n6911) );
  AN2HHD U9302 ( .I1(n12086), .I2(n13844), .O(n6913) );
  AN2HHD U9303 ( .I1(n8718), .I2(n8701), .O(n6914) );
  NR2CHD U9304 ( .I1(n9454), .I2(n12836), .O(n6917) );
  INVLHD U9305 ( .I(n12880), .O(n12808) );
  AN2HHD U9306 ( .I1(n9886), .I2(n12935), .O(n6918) );
  AN2EHD U9307 ( .I1(n13098), .I2(n11852), .O(n6919) );
  AN2HHD U9308 ( .I1(n9812), .I2(n8384), .O(n6920) );
  AN2HHD U9309 ( .I1(n8967), .I2(n8966), .O(n6923) );
  XOR2EHD U9310 ( .I1(_i_CLEFIA128_CON_T_x _14), .I2(DOUT_110), .O(n6924) );
  INVDHD U9311 ( .I(n7224), .O(n8345) );
  BUFNHD U9312 ( .I(n13288), .O(n13339) );
  AN2HHD U9313 ( .I1(n8132), .I2(_i_CLEFIA128_state_reg _1), .O(n6927) );
  AN3EHD U9314 ( .I1(n8797), .I2(_i_CLEFIA128_keyK _127), .I3(_i_CLEFIA128_keyL _127), .O(n6928) );
  XNR2KHD U9315 ( .I1(n11660), .I2(n7064), .O(n6931) );
  INVMHD U9316 ( .I(n9841), .O(n9840) );
  INVNHD U9317 ( .I(n11612), .O(n9568) );
  AN2HHD U9318 ( .I1(n9529), .I2(n12192), .O(n6932) );
  AN2HHD U9319 ( .I1(n14081), .I2(n9667), .O(n6933) );
  ND2HHD U9320 ( .I1(n12181), .I2(n14051), .O(n8997) );
  AN3EHD U9321 ( .I1(n13234), .I2(n13066), .I3(n8061), .O(n6935) );
  AN3EHD U9322 ( .I1(n9605), .I2(n8253), .I3(n7842), .O(n6936) );
  AN3EHD U9323 ( .I1(n9462), .I2(n14043), .I3(n10296), .O(n6937) );
  OR2EHD U9324 ( .I1(n8264), .I2(n13458), .O(n6939) );
  AN2EHD U9325 ( .I1(n13066), .I2(n8329), .O(n6940) );
  INVNHD U9326 ( .I(n11505), .O(n7674) );
  NR2EHD U9327 ( .I1(n8903), .I2(n7546), .O(n6941) );
  AN2EHD U9328 ( .I1(n7039), .I2(n8014), .O(n6943) );
  ND2DHD U9329 ( .I1(n11117), .I2(n12765), .O(n6945) );
  AN3EHD U9330 ( .I1(n12767), .I2(n8607), .I3(n7539), .O(n6946) );
  AN2EHD U9331 ( .I1(n7206), .I2(n12586), .O(n6948) );
  AN2HHD U9332 ( .I1(n11510), .I2(n12731), .O(n6949) );
  AN2EHD U9333 ( .I1(n11382), .I2(n8101), .O(n6952) );
  AN2EHD U9334 ( .I1(n9687), .I2(n12559), .O(n6954) );
  AN3HHD U9335 ( .I1(n6956), .I2(n6946), .I3(n12580), .O(n6955) );
  AN2EHD U9336 ( .I1(n7657), .I2(n7307), .O(n6956) );
  AN3EHD U9337 ( .I1(n12560), .I2(n12559), .I3(n7156), .O(n6957) );
  INVNHD U9338 ( .I(n8201), .O(n7384) );
  AN2EHD U9339 ( .I1(n7440), .I2(n13513), .O(n6958) );
  AN2HHD U9340 ( .I1(n8583), .I2(n12298), .O(n6959) );
  AN3EHD U9341 ( .I1(n8628), .I2(n12153), .I3(n13838), .O(n6961) );
  AN3EHD U9342 ( .I1(n13832), .I2(n9814), .I3(n8628), .O(n6963) );
  AN2HHD U9343 ( .I1(n13823), .I2(n8614), .O(n6964) );
  AN2EHD U9344 ( .I1(n13814), .I2(n13815), .O(n6965) );
  AN2HHD U9345 ( .I1(n10253), .I2(n10085), .O(n6966) );
  ND2KHD U9346 ( .I1(n7723), .I2(n10123), .O(n10960) );
  AN2EHD U9347 ( .I1(n10818), .I2(n12717), .O(n6967) );
  AN2HHD U9348 ( .I1(n8194), .I2(n10893), .O(n6969) );
  OR2KHD U9349 ( .I1(n9844), .I2(n10959), .O(n6970) );
  AN2EHD U9350 ( .I1(n10964), .I2(n10825), .O(n6971) );
  AN2EHD U9351 ( .I1(n12790), .I2(n7454), .O(n6972) );
  AN2HHD U9352 ( .I1(n8591), .I2(n12872), .O(n6973) );
  NR3BHD U9353 ( .I1(n12883), .I2(n12882), .I3(n12881), .O(n6974) );
  AN2EHD U9354 ( .I1(n7247), .I2(n10964), .O(n6976) );
  AN3EHD U9355 ( .I1(n8594), .I2(n6647), .I3(n8592), .O(n6977) );
  OR2HHD U9356 ( .I1(n7767), .I2(n8937), .O(n6978) );
  AN2EHD U9357 ( .I1(n9873), .I2(n9847), .O(n6979) );
  AN2EHD U9358 ( .I1(n9873), .I2(n13448), .O(n6980) );
  OR2EHD U9359 ( .I1(n8884), .I2(n9234), .O(n6981) );
  AN2EHD U9360 ( .I1(n13406), .I2(n6770), .O(n6982) );
  AN2HHD U9361 ( .I1(n12253), .I2(n13386), .O(n6985) );
  ND2KHD U9362 ( .I1(n7161), .I2(n7864), .O(n12635) );
  AN2EHD U9363 ( .I1(n10632), .I2(n10668), .O(n6988) );
  AN2HHD U9364 ( .I1(n7606), .I2(n12522), .O(n6989) );
  AN2EHD U9365 ( .I1(n11253), .I2(n7580), .O(n6990) );
  AN3HHD U9366 ( .I1(n7365), .I2(n12637), .I3(n11079), .O(n6993) );
  AN2EHD U9367 ( .I1(n12521), .I2(n6806), .O(n6995) );
  AN2EHD U9368 ( .I1(n7197), .I2(n7358), .O(n6996) );
  INVMHD U9369 ( .I(n9329), .O(n9042) );
  AN2HHD U9370 ( .I1(n9116), .I2(n9531), .O(n6998) );
  INVMHD U9371 ( .I(n10719), .O(n12456) );
  AN2HHD U9372 ( .I1(n9443), .I2(n11555), .O(n7000) );
  AN2HHD U9373 ( .I1(n11552), .I2(n11553), .O(n7001) );
  AN3HHD U9374 ( .I1(n12478), .I2(n11295), .I3(n12448), .O(n7002) );
  ND2KHD U9375 ( .I1(n8868), .I2(n9643), .O(n8031) );
  ND2HHD U9376 ( .I1(n12383), .I2(n12915), .O(n12280) );
  AN2HHD U9377 ( .I1(n9127), .I2(n13191), .O(n7007) );
  AN2EHD U9378 ( .I1(n9127), .I2(n13614), .O(n7009) );
  AN2EHD U9379 ( .I1(n12126), .I2(n13592), .O(n7011) );
  AN3EHD U9380 ( .I1(n12947), .I2(n7858), .I3(n12948), .O(n7012) );
  XNR2KHD U9381 ( .I1(n14367), .I2(n13938), .O(n15377) );
  ND3CHD U9382 ( .I1(n8613), .I2(n11765), .I3(n7353), .O(n9564) );
  BUFQHD U9383 ( .I(n12190), .O(n9186) );
  ND3CHD U9384 ( .I1(n12732), .I2(n12731), .I3(n7309), .O(n12733) );
  BUFKHD U9385 ( .I(n12449), .O(n9593) );
  ND2KHD U9386 ( .I1(n8524), .I2(n10071), .O(n8523) );
  ND3CHD U9387 ( .I1(n12585), .I2(n9625), .I3(n11323), .O(n11033) );
  ND2DHD U9388 ( .I1(n8011), .I2(n11130), .O(n9546) );
  INVGHD U9389 ( .I(n12504), .O(n10986) );
  ND2HHD U9390 ( .I1(n10437), .I2(n9581), .O(n9703) );
  BUFQHD U9391 ( .I(n10721), .O(n9903) );
  OA12HHD U9392 ( .B1(n13181), .B2(n12382), .A1(n13585), .O(n9602) );
  NR2EHD U9393 ( .I1(n10754), .I2(n10898), .O(n10757) );
  ND2KHD U9394 ( .I1(n10888), .I2(n12867), .O(n10898) );
  ND3CHD U9395 ( .I1(n10099), .I2(n9221), .I3(n13438), .O(n10098) );
  BUFQHD U9396 ( .I(n11907), .O(n12327) );
  ND3CHD U9397 ( .I1(n11219), .I2(n10374), .I3(n10373), .O(n10381) );
  ND2HHD U9398 ( .I1(n9811), .I2(n9807), .O(n7931) );
  ND2KHD U9399 ( .I1(n9916), .I2(n10825), .O(n12799) );
  ND2DHD U9400 ( .I1(n10453), .I2(n8233), .O(n8530) );
  BUFHHD U9401 ( .I(n12393), .O(n9752) );
  AN3EHD U9402 ( .I1(n12393), .I2(n12401), .I3(n10080), .O(n9520) );
  ND2HHD U9403 ( .I1(n13373), .I2(n9873), .O(n7268) );
  INVNHD U9404 ( .I(n10198), .O(n11614) );
  AN3B1HHD U9405 ( .I1(n10896), .I2(n9590), .B1(n8971), .O(n8548) );
  ND2HHD U9406 ( .I1(n12797), .I2(n12669), .O(n8918) );
  NR2EHD U9407 ( .I1(n13059), .I2(n13060), .O(n9630) );
  INVHHD U9408 ( .I(n11541), .O(n11551) );
  ND2DHD U9409 ( .I1(n12727), .I2(n11485), .O(n10517) );
  INVHHD U9410 ( .I(n14080), .O(n9507) );
  NR2CHD U9411 ( .I1(n7674), .I2(n11334), .O(n8537) );
  ND2DHD U9412 ( .I1(n15207), .I2(n15500), .O(n13969) );
  ND2DHD U9413 ( .I1(n13880), .I2(n13879), .O(n6101) );
  XNR2HHD U9414 ( .I1(n14489), .I2(n9757), .O(n14491) );
  ND2DHD U9415 ( .I1(n9535), .I2(n7860), .O(n10246) );
  INVDHD U9416 ( .I(n11201), .O(n11202) );
  ND3CHD U9417 ( .I1(n9365), .I2(n8336), .I3(n9375), .O(n9364) );
  ND2DHD U9418 ( .I1(n7020), .I2(n13421), .O(n9439) );
  INVGHD U9419 ( .I(n8084), .O(n7355) );
  INVGHD U9420 ( .I(n13422), .O(n7020) );
  INVHHD U9421 ( .I(n8004), .O(n7473) );
  INVCKGHD U9422 ( .I(n12385), .O(n12375) );
  BUFIHD U9423 ( .I(n11401), .O(n8863) );
  NR2EHD U9424 ( .I1(n7360), .I2(n11324), .O(n8013) );
  INVJHD U9425 ( .I(n10992), .O(n9231) );
  ND2DHD U9426 ( .I1(n14448), .I2(n14738), .O(n6366) );
  ND2DHD U9427 ( .I1(n14424), .I2(n14741), .O(n6373) );
  MUX2CHD U9428 ( .A(n14743), .B(n14742), .S(_i_CLEFIA128_CON_T_reg_4 ), .O(n14458) );
  MUX2CHD U9429 ( .A(n14743), .B(n14742), .S(_i_CLEFIA128_CON_T_xi _11), .O(n14453) );
  MUX2CHD U9430 ( .A(n14743), .B(n14742), .S(_i_CLEFIA128_CON_T_xi _9), .O(n14463) );
  INVKHD U9431 ( .I(n7384), .O(n8200) );
  BUFHHD U9432 ( .I(n8329), .O(n14087) );
  BUFLHD U9433 ( .I(n9208), .O(n7376) );
  OA12EHD U9434 ( .B1(n15499), .B2(n15224), .A1(n14105), .O(n14111) );
  OA12CHD U9435 ( .B1(n15499), .B2(n14814), .A1(n14165), .O(n14166) );
  OA12EHD U9436 ( .B1(n13277), .B2(n7143), .A1(n14922), .O(n8262) );
  OA12EHD U9437 ( .B1(n15499), .B2(n14383), .A1(n14341), .O(n8241) );
  OA12CHD U9438 ( .B1(n15499), .B2(n15393), .A1(n15068), .O(n8243) );
  OA12EHD U9439 ( .B1(n13277), .B2(n14927), .A1(n14835), .O(n14836) );
  OA12EHD U9440 ( .B1(n13277), .B2(n15280), .A1(n14963), .O(n8305) );
  OA12EHD U9441 ( .B1(n13277), .B2(n14923), .A1(n14840), .O(n14841) );
  OA12EHD U9442 ( .B1(n15499), .B2(n15316), .A1(n15308), .O(n8342) );
  OA12CHD U9443 ( .B1(n15499), .B2(n14802), .A1(n14801), .O(n8311) );
  OA12EHD U9444 ( .B1(n15499), .B2(n15488), .A1(n15487), .O(n15489) );
  OA12EHD U9445 ( .B1(n13277), .B2(n15125), .A1(n15093), .O(n15094) );
  OA12EHD U9446 ( .B1(n15499), .B2(n15330), .A1(n14642), .O(n14643) );
  OA12EHD U9447 ( .B1(n15499), .B2(n15345), .A1(n14270), .O(n14271) );
  OA12EHD U9448 ( .B1(n15499), .B2(n15141), .A1(n14571), .O(n14572) );
  OA12EHD U9449 ( .B1(n15499), .B2(n14608), .A1(n14607), .O(n14609) );
  OA12EHD U9450 ( .B1(n13277), .B2(n15073), .A1(n15072), .O(n8307) );
  OA12EHD U9451 ( .B1(n15499), .B2(n15159), .A1(n14807), .O(n14808) );
  OA12EHD U9452 ( .B1(n13277), .B2(n15306), .A1(n15305), .O(n8360) );
  OA12EHD U9453 ( .B1(n13277), .B2(n15074), .A1(n14992), .O(n8385) );
  OA12EHD U9454 ( .B1(n15499), .B2(n14866), .A1(n14010), .O(n8356) );
  AN2EHD U9455 ( .I1(n14468), .I2(n14725), .O(n14473) );
  OA12EHD U9456 ( .B1(n15499), .B2(n14924), .A1(n12446), .O(n12447) );
  ND2DHD U9457 ( .I1(n14718), .I2(n14717), .O(n6367) );
  OA12EHD U9458 ( .B1(n13277), .B2(n15415), .A1(n15138), .O(n15139) );
  OA12EHD U9459 ( .B1(n13277), .B2(n15249), .A1(n15248), .O(n15250) );
  ND2DHD U9460 ( .I1(n14408), .I2(n14741), .O(n6374) );
  NR2CHD U9461 ( .I1(n14411), .I2(n14716), .O(n14417) );
  NR2IHD U9462 ( .I1(n14444), .I2(n14475), .O(n14433) );
  OA112CHD U9463 ( .C1(n15422), .C2(n15189), .A1(n15188), .B1(n15187), .O(n15190) );
  NR2IHD U9464 ( .I1(n14434), .I2(n14752), .O(n14465) );
  AN2CHD U9465 ( .I1(n15253), .I2(n9501), .O(n15256) );
  INVNHD U9466 ( .I(n8177), .O(n8178) );
  OA112EHD U9467 ( .C1(n14383), .C2(n15513), .A1(n10934), .B1(n10933), .O(n8328) );
  NR2CHD U9468 ( .I1(n10926), .I2(n10925), .O(n10927) );
  AN2CHD U9469 ( .I1(n15252), .I2(n8448), .O(n9501) );
  INVLHD U9470 ( .I(n9744), .O(n10939) );
  NR2CHD U9471 ( .I1(n15319), .I2(n15318), .O(n15320) );
  AN2HHD U9472 ( .I1(n11727), .I2(n11721), .O(n13835) );
  AN2CHD U9473 ( .I1(n13275), .I2(n13274), .O(n13276) );
  AN2HHD U9474 ( .I1(n11736), .I2(n11721), .O(n13826) );
  NR2BHD U9475 ( .I1(n9500), .I2(n9499), .O(n14854) );
  INVJHD U9476 ( .I(n7360), .O(n11378) );
  INVJHD U9477 ( .I(n14432), .O(n14475) );
  NR2CHD U9478 ( .I1(n14396), .I2(n14395), .O(n14397) );
  BUFQHD U9479 ( .I(n14796), .O(n15422) );
  NR2CHD U9480 ( .I1(n14323), .I2(n14322), .O(n14324) );
  AN2HHD U9481 ( .I1(n12054), .I2(n12053), .O(n13585) );
  INVDHD U9482 ( .I(n14713), .O(n14420) );
  INVGHD U9483 ( .I(n10938), .O(n9020) );
  INVCHD U9484 ( .I(n11130), .O(n7603) );
  INVQHD U9485 ( .I(n15416), .O(n7043) );
  INVIHD U9486 ( .I(n9591), .O(n10690) );
  BUFLHD U9487 ( .I(n11129), .O(n15512) );
  INVNHD U9488 ( .I(n11129), .O(n11130) );
  XNR2HHD U9489 ( .I1(n10610), .I2(n10609), .O(n11318) );
  INVDHD U9490 ( .I(n14407), .O(n14404) );
  INVQHD U9491 ( .I(n15513), .O(n15500) );
  AOI22BHD U9492 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _100), .B1(n15504), .B2(_i_CLEFIA128_keyK _36), .O(n13265) );
  AO22CHD U9493 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _68), .B1(n15504), .B2(_i_CLEFIA128_keyK _4), .O(n8390) );
  AO22CHD U9494 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _75), .B1(n15504), .B2(_i_CLEFIA128_keyK _11), .O(n15321) );
  AO22CHD U9495 ( .A1(n7045), .A2(n15310), .B1(n15504), .B2(n15309), .O(n15311) );
  INVMHD U9496 ( .I(n7866), .O(n7016) );
  AO22CHD U9497 ( .A1(n7045), .A2(n13985), .B1(n15504), .B2(n13984), .O(n13986) );
  AOI22BHD U9498 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _106), .B1(n15504), .B2(_i_CLEFIA128_keyK _42), .O(n14353) );
  AO22CHD U9499 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _66), .B1(n15504), .B2(_i_CLEFIA128_keyK _2), .O(n13927) );
  AO22CHD U9500 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _94), .B1(n15504), .B2(_i_CLEFIA128_keyK _30), .O(n13913) );
  AO22CHD U9501 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _102), .B1(n15504), .B2(_i_CLEFIA128_keyK _38), .O(n13852) );
  INVDHD U9502 ( .I(n10912), .O(n14435) );
  NR2EHD U9503 ( .I1(SRST), .I2(n14402), .O(n14407) );
  NR2GHD U9504 ( .I1(n14444), .I2(n8627), .O(n14427) );
  INVMHD U9505 ( .I(n10300), .O(n7045) );
  NR2BHD U9506 ( .I1(n15014), .I2(n13277), .O(n14640) );
  NR2CHD U9507 ( .I1(n8626), .I2(n7103), .O(n12011) );
  ND2HHD U9508 ( .I1(n13280), .I2(n13279), .O(n13281) );
  INVNHD U9509 ( .I(n8222), .O(n15504) );
  AN2EHD U9510 ( .I1(n14399), .I2(n14683), .O(n14723) );
  NR2CHD U9511 ( .I1(n14415), .I2(n6741), .O(n13283) );
  ND2KHD U9512 ( .I1(n15492), .I2(n10911), .O(n10912) );
  INVQHD U9513 ( .I(n13292), .O(n13277) );
  OR2EHD U9514 ( .I1(n14400), .I2(n13292), .O(n14401) );
  ND2DHD U9515 ( .I1(n7389), .I2(n6928), .O(n8132) );
  ND2KHD U9516 ( .I1(n14688), .I2(n10302), .O(n8222) );
  BUFNHD U9517 ( .I(n12895), .O(n15492) );
  ND2HHD U9518 ( .I1(n11879), .I2(_i_CLEFIA128_keyL _105), .O(n11878) );
  NR2CHD U9519 ( .I1(n14678), .I2(n14719), .O(n13284) );
  NR2EHD U9520 ( .I1(n13286), .I2(n14685), .O(n13291) );
  NR2EHD U9521 ( .I1(n11862), .I2(n8439), .O(n8124) );
  INVNHD U9522 ( .I(n8259), .O(n7017) );
  INVDHD U9523 ( .I(_i_CLEFIA128_keyL _63), .O(n15421) );
  INVDHD U9524 ( .I(_i_CLEFIA128_keyL _23), .O(n15040) );
  INVDHD U9525 ( .I(_i_CLEFIA128_keyL _108), .O(n15349) );
  INVDHD U9526 ( .I(_i_CLEFIA128_keyL _127), .O(n15423) );
  INVDHD U9527 ( .I(_i_CLEFIA128_keyL _44), .O(n15042) );
  INVCHD U9528 ( .I(_i_CLEFIA128_keyL _110), .O(n7392) );
  INVDHD U9529 ( .I(DOUT_120), .O(n14608) );
  INVDHD U9530 ( .I(_i_CLEFIA128_keyL _96), .O(n14945) );
  INVMHD U9531 ( .I(_i_CLEFIA128_keyL _26), .O(n15277) );
  XNR2EHD U9532 ( .I1(_i_CLEFIA128_CON_T_xi _13), .I2(DOUT_111), .O(n8404));
  INVDHD U9533 ( .I(_i_CLEFIA128_keyL _62), .O(n15100) );
  INVDHD U9534 ( .I(_i_CLEFIA128_keyL _126), .O(n15233) );
  INVDHD U9535 ( .I(_i_CLEFIA128_keyL _119), .O(n15239) );
  INVDHD U9536 ( .I(_i_CLEFIA128_keyL _55), .O(n15121) );
  XNR2EHD U9537 ( .I1(_i_CLEFIA128_CON_T_x _8), .I2(DOUT_119), .O(n11695) );
  INVDHD U9538 ( .I(_i_CLEFIA128_keyL _122), .O(n15341) );
  INVDHD U9539 ( .I(_i_CLEFIA128_keyL _2), .O(n15029) );
  INVDHD U9540 ( .I(_i_CLEFIA128_keyL _115), .O(n15348) );
  INVDHD U9541 ( .I(_i_CLEFIA128_keyL _114), .O(n15205) );
  INVDHD U9542 ( .I(_i_CLEFIA128_keyL _97), .O(n15284) );
  XNR2EHD U9543 ( .I1(_i_CLEFIA128_CON_T_x _7), .I2(DOUT_54), .O(n10582) );
  INVDHD U9544 ( .I(_i_CLEFIA128_keyL _47), .O(n15289) );
  INVMHD U9545 ( .I(_i_CLEFIA128_keyL _35), .O(n15058) );
  INVDHD U9546 ( .I(_i_CLEFIA128_keyL _54), .O(n15290) );
  INVDHD U9547 ( .I(_i_CLEFIA128_keyL _111), .O(n15267) );
  INVDHD U9548 ( .I(_i_CLEFIA128_keyL _118), .O(n15254) );
  INVJHD U9549 ( .I(_i_CLEFIA128_keyK _80), .O(n13778) );
  INVDHD U9550 ( .I(_i_CLEFIA128_keyL _121), .O(n15214) );
  INVKHD U9551 ( .I(_i_CLEFIA128_state_reg _0), .O(n10301) );
  INVMHD U9552 ( .I(_i_CLEFIA128_keyL _33), .O(n15280) );
  INVKHD U9553 ( .I(_i_CLEFIA128_keyL _32), .O(n14954) );
  NR2BHD U9554 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(_i_CLEFIA128_keyK _118), .O(n11696) );
  NR2CHD U9555 ( .I1(_i_CLEFIA128_rndcnt_reg _2), .I2(_i_CLEFIA128_rndcnt_reg _4), .O(n13282) );
  XNR2EHD U9556 ( .I1(_i_CLEFIA128_CON_T_x _7), .I2(DOUT_103), .O(n12014) );
  INVCHD U9557 ( .I(DOUT_29), .O(n7073) );
  INVCHD U9558 ( .I(DOUT_93), .O(n7956) );
  INVCHD U9559 ( .I(_i_CLEFIA128_keyL _48), .O(n15125) );
  INVDHD U9560 ( .I(DOUT_88), .O(n9408) );
  INVCHD U9561 ( .I(DOUT_70), .O(n8064) );
  INVDHD U9562 ( .I(DOUT_56), .O(n14880) );
  ND2KHD U9563 ( .I1(_i_CLEFIA128_state_reg _1), .I2(_i_CLEFIA128_state_reg _0), .O(n14444) );
  INVDHD U9564 ( .I(_i_CLEFIA128_keyL _100), .O(n15169) );
  INVDHD U9565 ( .I(_i_CLEFIA128_rndcnt_reg _2), .O(n14412) );
  INVCHD U9566 ( .I(_i_CLEFIA128_keyK _0), .O(n8777) );
  ND2CHD U9567 ( .I1(_i_CLEFIA128_keyK _6), .I2(_i_CLEFIA128_keyL _6), .O(n9472) );
  INVDHD U9568 ( .I(DOUT_113), .O(n14871) );
  INVCHD U9569 ( .I(DOUT_84), .O(n10181) );
  INVKHD U9570 ( .I(_i_CLEFIA128_keyL _113), .O(n8662) );
  INVDHD U9571 ( .I(_i_CLEFIA128_keyL _38), .O(n14976) );
  INVDHD U9572 ( .I(_i_CLEFIA128_keyL _102), .O(n14557) );
  INVDHD U9573 ( .I(_i_CLEFIA128_keyL _31), .O(n14975) );
  INVKHD U9574 ( .I(_i_CLEFIA128_keyL _28), .O(n15298) );
  INVMHD U9575 ( .I(KEYSET), .O(n10913) );
  ND3CHD U9576 ( .I1(n10197), .I2(n7604), .I3(n10927), .O(n6123) );
  ND3CHD U9577 ( .I1(n7211), .I2(n7210), .I3(n15013), .O(n6167) );
  ND2DHD U9578 ( .I1(n8730), .I2(n14632), .O(n6273) );
  ND2DHD U9579 ( .I1(n7352), .I2(n15094), .O(n6272) );
  ND2HHD U9580 ( .I1(n15486), .I2(n14774), .O(n14782) );
  ND2DHD U9581 ( .I1(n9147), .I2(n14530), .O(n6334) );
  INVJHD U9582 ( .I(n9010), .O(n14168) );
  ND2HHD U9583 ( .I1(n13112), .I2(n13111), .O(n12949) );
  OA12EHD U9584 ( .B1(n9071), .B2(n12083), .A1(n13817), .O(n12084) );
  INVGHD U9585 ( .I(n13467), .O(n9254) );
  INVIHD U9586 ( .I(n13064), .O(n13493) );
  NR2EHD U9587 ( .I1(n12884), .I2(n8580), .O(n7740) );
  ND2DHD U9588 ( .I1(n8249), .I2(n11557), .O(n9798) );
  NR2EHD U9589 ( .I1(n9347), .I2(n9346), .O(n9345) );
  INVJHD U9590 ( .I(n12532), .O(n7018) );
  ND3CHD U9591 ( .I1(n13092), .I2(n13093), .I3(n13091), .O(n13094) );
  NR2GHD U9592 ( .I1(n7690), .I2(n7689), .O(n7688) );
  NR2EHD U9593 ( .I1(n13525), .I2(n13524), .O(n13527) );
  NR2EHD U9594 ( .I1(n7461), .I2(n7459), .O(n7462) );
  ND2DHD U9595 ( .I1(n8996), .I2(n9230), .O(n12182) );
  AN3EHD U9596 ( .I1(n14047), .I2(n8667), .I3(n9230), .O(n8666) );
  ND2HHD U9597 ( .I1(n8086), .I2(n9814), .O(n13547) );
  INVJHD U9598 ( .I(n12634), .O(n10171) );
  NR2EHD U9599 ( .I1(n7279), .I2(n12572), .O(n7278) );
  ND2HHD U9600 ( .I1(n8921), .I2(n9590), .O(n7733) );
  NR2EHD U9601 ( .I1(n12991), .I2(n9928), .O(n9927) );
  NR2GHD U9602 ( .I1(n11140), .I2(n11139), .O(n11147) );
  NR2EHD U9603 ( .I1(n13197), .I2(n13196), .O(n13204) );
  INVCKIHD U9604 ( .I(n11305), .O(n11308) );
  ND2HHD U9605 ( .I1(n9310), .I2(n12868), .O(n7889) );
  NR2EHD U9606 ( .I1(n8419), .I2(n9015), .O(n10294) );
  INVLHD U9607 ( .I(n9436), .O(n13421) );
  NR2EHD U9608 ( .I1(n8609), .I2(n7264), .O(n8608) );
  NR2EHD U9609 ( .I1(n9653), .I2(n12002), .O(n12003) );
  ND2DHD U9610 ( .I1(n13630), .I2(n7552), .O(n13632) );
  INVGHD U9611 ( .I(n11062), .O(n7194) );
  NR2EHD U9612 ( .I1(n10705), .I2(n11139), .O(n10706) );
  NR2EHD U9613 ( .I1(n12587), .I2(n12588), .O(n9025) );
  INVJHD U9614 ( .I(n12720), .O(n9619) );
  INVIHD U9615 ( .I(n8965), .O(n7022) );
  NR2GHD U9616 ( .I1(n10285), .I2(n7891), .O(n7884) );
  INVJHD U9617 ( .I(n13088), .O(n13473) );
  INVKHD U9618 ( .I(n12621), .O(n7024) );
  INVGHD U9619 ( .I(n9648), .O(n10077) );
  INVKHD U9620 ( .I(n12757), .O(n7025) );
  NR2EHD U9621 ( .I1(n10762), .I2(n6767), .O(n9385) );
  INVIHD U9622 ( .I(n9575), .O(n10673) );
  AN2CHD U9623 ( .I1(n14743), .I2(n14440), .O(n14442) );
  BUFGHD U9624 ( .I(n8215), .O(n10889) );
  ND2DHD U9625 ( .I1(n11026), .I2(n7498), .O(n11027) );
  ND2DHD U9626 ( .I1(n8247), .I2(n7306), .O(n10539) );
  BUFCKEHD U9627 ( .I(n13671), .O(n9098) );
  ND2DHD U9628 ( .I1(n14061), .I2(n14062), .O(n9182) );
  ND3CHD U9629 ( .I1(n8581), .I2(n13844), .I3(n13810), .O(n11726) );
  ND2CHD U9630 ( .I1(n14433), .I2(_i_CLEFIA128_CON_T_x _7), .O(n14734) );
  ND2CHD U9631 ( .I1(n14433), .I2(_i_CLEFIA128_CON_T_x _9), .O(n14729) );
  INVGHD U9632 ( .I(n10069), .O(n7028) );
  ND2KHD U9633 ( .I1(n9183), .I2(n9184), .O(n14063) );
  AO222CHD U9634 ( .A1(n14475), .A2(_i_CLEFIA128_CON_T_x _7), .B1(n14465), .B2(_i_CLEFIA128_CON_T_x _8), .C1(_i_CLEFIA128_CON_T_x _6), .C2(n14433), .O(n6359) );
  AN2EHD U9635 ( .I1(n11403), .I2(n12564), .O(n11404) );
  NR2CHD U9636 ( .I1(n14554), .I2(n14553), .O(n14555) );
  NR2CHD U9637 ( .I1(n14599), .I2(n14598), .O(n14600) );
  NR2CHD U9638 ( .I1(n14497), .I2(n14496), .O(n14498) );
  OA12CHD U9639 ( .B1(n15499), .B2(n15483), .A1(n15482), .O(n15484) );
  NR2CHD U9640 ( .I1(n14523), .I2(n14522), .O(n14524) );
  NR2CHD U9641 ( .I1(n14487), .I2(n14486), .O(n14488) );
  NR2CHD U9642 ( .I1(n14503), .I2(n14502), .O(n14504) );
  NR2CHD U9643 ( .I1(n14534), .I2(n14533), .O(n14535) );
  NR2CHD U9644 ( .I1(n14662), .I2(n14661), .O(n14663) );
  NR2CHD U9645 ( .I1(n14652), .I2(n14651), .O(n14653) );
  NR2CHD U9646 ( .I1(n14631), .I2(n14630), .O(n14632) );
  NR2CHD U9647 ( .I1(n14594), .I2(n14593), .O(n14595) );
  AN2CHD U9648 ( .I1(n14865), .I2(n8449), .O(n8255) );
  NR2CHD U9649 ( .I1(n14569), .I2(n14568), .O(n14570) );
  ND2CHD U9650 ( .I1(n9184), .I2(n14060), .O(n8331) );
  NR2CHD U9651 ( .I1(n14549), .I2(n14548), .O(n14550) );
  NR2CHD U9652 ( .I1(n14589), .I2(n14588), .O(n14590) );
  NR2CHD U9653 ( .I1(n14518), .I2(n14517), .O(n14519) );
  ND2DHD U9654 ( .I1(n14465), .I2(n14464), .O(n14737) );
  OA12CHD U9655 ( .B1(n15499), .B2(n15491), .A1(n15490), .O(n8281) );
  BUFIHD U9656 ( .I(n14044), .O(n9529) );
  NR2CHD U9657 ( .I1(n14584), .I2(n14583), .O(n14585) );
  NR2CHD U9658 ( .I1(n14625), .I2(n14624), .O(n14626) );
  NR2CHD U9659 ( .I1(n14667), .I2(n14666), .O(n14668) );
  AN2CHD U9660 ( .I1(n14468), .I2(n14460), .O(n14462) );
  NR2CHD U9661 ( .I1(n14619), .I2(n14618), .O(n14620) );
  NR2CHD U9662 ( .I1(n14579), .I2(n14578), .O(n14580) );
  NR2CHD U9663 ( .I1(n14561), .I2(n14560), .O(n14562) );
  NR2CHD U9664 ( .I1(n14513), .I2(n14512), .O(n14514) );
  NR2CHD U9665 ( .I1(n14640), .I2(n14639), .O(n14641) );
  BUFQHD U9666 ( .I(n11892), .O(n7032) );
  NR2CHD U9667 ( .I1(n14539), .I2(n14538), .O(n14540) );
  NR2CHD U9668 ( .I1(n14605), .I2(n14604), .O(n14606) );
  INVJHD U9669 ( .I(n12809), .O(n7033) );
  OA12CHD U9670 ( .B1(n15499), .B2(n15386), .A1(n13861), .O(n13863) );
  NR2CHD U9671 ( .I1(n14508), .I2(n14507), .O(n14509) );
  NR2CHD U9672 ( .I1(n14481), .I2(n14480), .O(n14482) );
  OA12CHD U9673 ( .B1(n15499), .B2(n15511), .A1(n13748), .O(n13749) );
  NR2CHD U9674 ( .I1(n14544), .I2(n14543), .O(n14545) );
  AO12CHD U9675 ( .B1(n14716), .B2(n14715), .A1(n14714), .O(n6371) );
  NR2BHD U9676 ( .I1(n14714), .I2(n14418), .O(n14416) );
  OA112CHD U9677 ( .C1(n15422), .C2(n15092), .A1(n15091), .B1(n15090), .O(n15093) );
  INVNHD U9678 ( .I(n8292), .O(n7035) );
  OA112CHD U9679 ( .C1(n15422), .C2(n14864), .A1(n14863), .B1(n14862), .O(n14865) );
  OA112CHD U9680 ( .C1(n15290), .C2(n15420), .A1(n14855), .B1(n14854), .O(n14857) );
  OA112CHD U9681 ( .C1(n15422), .C2(n15186), .A1(n14897), .B1(n14896), .O(n14898) );
  ND2DHD U9682 ( .I1(n7904), .I2(n7720), .O(n8371) );
  OA112CHD U9683 ( .C1(n15422), .C2(n15270), .A1(n14962), .B1(n14961), .O(n14963) );
  INVNHD U9684 ( .I(n12141), .O(n15499) );
  OA112CHD U9685 ( .C1(n15422), .C2(n15050), .A1(n15038), .B1(n15037), .O(n15039) );
  OA112CHD U9686 ( .C1(n15422), .C2(n15185), .A1(n15174), .B1(n15173), .O(n15175) );
  OA112CHD U9687 ( .C1(n15422), .C2(n15036), .A1(n14798), .B1(n14797), .O(n14799) );
  OA112CHD U9688 ( .C1(n15422), .C2(n15201), .A1(n14810), .B1(n14809), .O(n14811) );
  AO12CHD U9689 ( .B1(BSY), .B2(n14726), .A1(n14748), .O(n6503) );
  OA112CHD U9690 ( .C1(n15422), .C2(n15426), .A1(n15411), .B1(n15410), .O(n15412) );
  OA112CHD U9691 ( .C1(n15422), .C2(n14918), .A1(n14910), .B1(n14909), .O(n14911) );
  OA112CHD U9692 ( .C1(n15422), .C2(n15296), .A1(n15295), .B1(n15294), .O(n15297) );
  INVCHD U9693 ( .I(n13458), .O(n13413) );
  AN2CHD U9694 ( .I1(n14741), .I2(n14455), .O(n14457) );
  AN2CHD U9695 ( .I1(n14741), .I2(n14450), .O(n14452) );
  ND2CHD U9696 ( .I1(n14741), .I2(n14740), .O(n14744) );
  ND2DHD U9697 ( .I1(n14748), .I2(n14435), .O(n14468) );
  OA112CHD U9698 ( .C1(n15422), .C2(n15301), .A1(n15071), .B1(n15070), .O(n15072) );
  OA112CHD U9699 ( .C1(n15422), .C2(n14930), .A1(n14921), .B1(n14920), .O(n14922) );
  NR2CHD U9700 ( .I1(n14038), .I2(n14037), .O(n14039) );
  NR2CHD U9701 ( .I1(n14780), .I2(n14779), .O(n14781) );
  NR2CHD U9702 ( .I1(n14293), .I2(n14292), .O(n14294) );
  OR2CHD U9703 ( .I1(n14449), .I2(n14432), .O(n14450) );
  NR2BHD U9704 ( .I1(n14727), .I2(n14432), .O(n14728) );
  NR2CHD U9705 ( .I1(n15008), .I2(n15007), .O(n15009) );
  NR2CHD U9706 ( .I1(n14024), .I2(n14023), .O(n14025) );
  NR2CHD U9707 ( .I1(n13878), .I2(n13877), .O(n13879) );
  NR2CHD U9708 ( .I1(n15226), .I2(n15225), .O(n15227) );
  NR2CHD U9709 ( .I1(n14238), .I2(n14237), .O(n14239) );
  NR2CHD U9710 ( .I1(n14892), .I2(n14891), .O(n14893) );
  OA112CHD U9711 ( .C1(n15423), .C2(n15420), .A1(n13357), .B1(n13356), .O(n13359) );
  NR2CHD U9712 ( .I1(n14702), .I2(n14701), .O(n14703) );
  NR2CHD U9713 ( .I1(n14002), .I2(n14001), .O(n14003) );
  OA112CHD U9714 ( .C1(n7143), .C2(n15420), .A1(n14830), .B1(n14829), .O(n14832) );
  OR2CHD U9715 ( .I1(n14459), .I2(n14432), .O(n14460) );
  OA112CHD U9716 ( .C1(n15289), .C2(n15420), .A1(n15288), .B1(n15287), .O(n15292) );
  NR2CHD U9717 ( .I1(n14304), .I2(n14303), .O(n14305) );
  NR2CHD U9718 ( .I1(n14762), .I2(n14761), .O(n14763) );
  OA112CHD U9719 ( .C1(n15341), .C2(n15420), .A1(n15026), .B1(n15025), .O(n15028) );
  OA112CHD U9720 ( .C1(n15046), .C2(n15420), .A1(n15045), .B1(n15044), .O(n15049) );
  AN2HHD U9721 ( .I1(n12140), .I2(n15450), .O(n12141) );
  NR2CHD U9722 ( .I1(n14339), .I2(n14338), .O(n14340) );
  NR2CHD U9723 ( .I1(n14792), .I2(n14791), .O(n14793) );
  OA112CHD U9724 ( .C1(n15348), .C2(n15420), .A1(n15347), .B1(n15346), .O(n15351) );
  NR2CHD U9725 ( .I1(n14099), .I2(n14098), .O(n14100) );
  OR2CHD U9726 ( .I1(n14464), .I2(n14432), .O(n14440) );
  OA112CHD U9727 ( .C1(n15249), .C2(n15420), .A1(n15108), .B1(n15107), .O(n15110) );
  NR2CHD U9728 ( .I1(n15363), .I2(n15362), .O(n15364) );
  NR2CHD U9729 ( .I1(n13775), .I2(n13774), .O(n13776) );
  INVNHD U9730 ( .I(n8759), .O(n11176) );
  OA112CHD U9731 ( .C1(n15239), .C2(n15420), .A1(n15238), .B1(n15237), .O(n15241) );
  OR2CHD U9732 ( .I1(n14739), .I2(n14432), .O(n14740) );
  OA112CHD U9733 ( .C1(n15420), .C2(n14943), .A1(n14843), .B1(n14842), .O(n14845) );
  NR2CHD U9734 ( .I1(n13710), .I2(n13709), .O(n13711) );
  OR2CHD U9735 ( .I1(n14454), .I2(n14432), .O(n14455) );
  NR2CHD U9736 ( .I1(n13697), .I2(n13696), .O(n13698) );
  OA112CHD U9737 ( .C1(n14975), .C2(n15420), .A1(n14974), .B1(n14973), .O(n14978) );
  OA112CHD U9738 ( .C1(n14483), .C2(n15420), .A1(n13333), .B1(n13332), .O(n13335) );
  NR2CHD U9739 ( .I1(n13959), .I2(n13958), .O(n13960) );
  OA112CHD U9740 ( .C1(n14976), .C2(n15420), .A1(n14969), .B1(n14968), .O(n14971) );
  NR2CHD U9741 ( .I1(n14264), .I2(n14263), .O(n14265) );
  OA112CHD U9742 ( .C1(n15420), .C2(n15042), .A1(n13317), .B1(n13316), .O(n13319) );
  NR2CHD U9743 ( .I1(n15332), .I2(n15331), .O(n15333) );
  NR2CHD U9744 ( .I1(n15388), .I2(n15387), .O(n15389) );
  OA112CHD U9745 ( .C1(n7392), .C2(n15420), .A1(n14947), .B1(n14946), .O(n14949) );
  OA112CHD U9746 ( .C1(n15420), .C2(n15236), .A1(n15112), .B1(n15111), .O(n15114) );
  OA112CHD U9747 ( .C1(n15100), .C2(n15420), .A1(n15082), .B1(n15081), .O(n15084) );
  NR2CHD U9748 ( .I1(n14123), .I2(n14122), .O(n14124) );
  OA112CHD U9749 ( .C1(n15415), .C2(n15420), .A1(n14873), .B1(n14872), .O(n14875) );
  NR2CHD U9750 ( .I1(n13981), .I2(n13980), .O(n13982) );
  NR2CHD U9751 ( .I1(n14282), .I2(n14281), .O(n14283) );
  OA112CHD U9752 ( .C1(n15274), .C2(n15420), .A1(n15273), .B1(n15272), .O(n15276) );
  OR2EHD U9753 ( .I1(n12893), .I2(n12892), .O(n12894) );
  NR2CHD U9754 ( .I1(n14386), .I2(n14385), .O(n14387) );
  OA112CHD U9755 ( .C1(n15254), .C2(n15420), .A1(n14859), .B1(n14858), .O(n14861) );
  NR2CHD U9756 ( .I1(n15516), .I2(n15515), .O(n15517) );
  ND2HHD U9757 ( .I1(n14432), .I2(n14444), .O(n14752) );
  NR2CHD U9758 ( .I1(n14163), .I2(n14162), .O(n14164) );
  NR2CHD U9759 ( .I1(n14359), .I2(n14358), .O(n14360) );
  NR2CHD U9760 ( .I1(n14191), .I2(n14190), .O(n14192) );
  NR2CHD U9761 ( .I1(n13262), .I2(n13261), .O(n13263) );
  BUFQHD U9762 ( .I(n11942), .O(n7038) );
  NR2CHD U9763 ( .I1(n14374), .I2(n14373), .O(n14375) );
  OA112CHD U9764 ( .C1(n15403), .C2(n15420), .A1(n15402), .B1(n15401), .O(n15406) );
  NR2CHD U9765 ( .I1(n15464), .I2(n15463), .O(n15465) );
  OA112CHD U9766 ( .C1(n15214), .C2(n15420), .A1(n13313), .B1(n13312), .O(n13315) );
  BUFQHD U9767 ( .I(n10512), .O(n7039) );
  INVQHD U9768 ( .I(n8179), .O(n7040) );
  AN2EHD U9769 ( .I1(n15512), .I2(n12139), .O(n12140) );
  INVKHD U9770 ( .I(n8206), .O(n8205) );
  OA22CHD U9771 ( .A1(n15385), .A2(n15416), .B1(n13339), .B2(n15289), .O(n15278) );
  NR2BHD U9772 ( .I1(n15159), .I2(n15416), .O(n9500) );
  AN2HHD U9773 ( .I1(n12864), .I2(n12846), .O(n12671) );
  NR2CHD U9774 ( .I1(n14413), .I2(n14709), .O(n14714) );
  AN3CHD U9775 ( .I1(n14723), .I2(n15522), .I3(n14722), .O(n14726) );
  OR2CHD U9776 ( .I1(n9502), .I2(n15420), .O(n8448) );
  OA22CHD U9777 ( .A1(n14945), .A2(n15420), .B1(n14919), .B2(n13339), .O(n14910) );
  INVCHD U9778 ( .I(n14694), .O(n14691) );
  NR2BHD U9779 ( .I1(n9502), .I2(n13339), .O(n9499) );
  NR2BHD U9780 ( .I1(n15239), .I2(n13277), .O(n14605) );
  OA112CHD U9781 ( .C1(n10912), .C2(n10932), .A1(n10931), .B1(n10930), .O(n10934) );
  NR2BHD U9782 ( .I1(n15423), .I2(n13277), .O(n14529) );
  BUFNHD U9783 ( .I(n13281), .O(n15420) );
  NR2BHD U9784 ( .I1(n14690), .I2(n14689), .O(n14694) );
  ND2CHD U9785 ( .I1(n10928), .I2(DOUT_20), .O(n10931) );
  OR3CHD U9786 ( .I1(_i_CLEFIA128_keyK _122), .I2(n14678), .I3(n14683), .O(n14682) );
  ND2DHD U9787 ( .I1(n10501), .I2(n9474), .O(n9473) );
  OR2CHD U9788 ( .I1(n14412), .I2(n6722), .O(n14414) );
  NR2BHD U9789 ( .I1(n14684), .I2(n14683), .O(n14690) );
  OR2CHD U9790 ( .I1(n8222), .I2(n14483), .O(n14989) );
  NR2GHD U9791 ( .I1(n13292), .I2(n13291), .O(n13293) );
  AN2CHD U9792 ( .I1(n14688), .I2(n14687), .O(n14689) );
  OA12EHD U9793 ( .B1(n11604), .B2(_i_CLEFIA128_keyL _126), .A1(_i_CLEFIA128_state_reg _1), .O(n8152) );
  ND2DHD U9794 ( .I1(n11924), .I2(_i_CLEFIA128_keyL _47), .O(n7063) );
  OA12EHD U9795 ( .B1(n11922), .B2(_i_CLEFIA128_keyL _111), .A1(_i_CLEFIA128_state_reg _1), .O(n7388) );
  OA12EHD U9796 ( .B1(n11916), .B2(_i_CLEFIA128_keyL _110), .A1(_i_CLEFIA128_state_reg _1), .O(n7391) );
  ND2DHD U9797 ( .I1(n11918), .I2(_i_CLEFIA128_keyL _46), .O(n7145) );
  INVDHD U9798 ( .I(n14425), .O(n12139) );
  OA12EHD U9799 ( .B1(n8130), .B2(n7532), .A1(_i_CLEFIA128_state_reg _1), .O(n7531) );
  ND2HHD U9800 ( .I1(n10457), .I2(_i_CLEFIA128_state_reg _1), .O(n7482) );
  XNR2HHD U9801 ( .I1(_i_CLEFIA128_keyL _66), .I2(n7576), .O(n10470) );
  INVCHD U9802 ( .I(n14685), .O(n14680) );
  ND2HHD U9803 ( .I1(n8259), .I2(n10917), .O(n14425) );
  ND2HHD U9804 ( .I1(n7453), .I2(_i_CLEFIA128_state_reg _1), .O(n9771) );
  NR2BHD U9805 ( .I1(n14686), .I2(n14685), .O(n14687) );
  INVCHD U9806 ( .I(n14719), .O(n14720) );
  ND2CHD U9807 ( .I1(n13949), .I2(_i_CLEFIA128_rndcnt_reg _0), .O(n10392) );
  INVGHD U9808 ( .I(n11886), .O(n7812) );
  ND2HHD U9809 ( .I1(n8039), .I2(_i_CLEFIA128_keyK _56), .O(n7983) );
  ND2HHD U9810 ( .I1(n7219), .I2(_i_CLEFIA128_keyK _25), .O(n8038) );
  ND2CHD U9811 ( .I1(n13995), .I2(_i_CLEFIA128_rndcnt_reg _0), .O(n11699) );
  ND2CHD U9812 ( .I1(n10337), .I2(n13802), .O(n12018) );
  ND2CHD U9813 ( .I1(n14026), .I2(_i_CLEFIA128_rndcnt_reg _0), .O(n11917) );
  ND2CHD U9814 ( .I1(n8626), .I2(n9173), .O(n12010) );
  ND2CHD U9815 ( .I1(n13984), .I2(_i_CLEFIA128_rndcnt_reg _0), .O(n10576) );
  INVCHD U9816 ( .I(n14434), .O(n14400) );
  AN2EHD U9817 ( .I1(n7220), .I2(n8798), .O(n10298) );
  ND2CHD U9818 ( .I1(n13765), .I2(_i_CLEFIA128_rndcnt_reg _0), .O(n11689) );
  NR2BHD U9819 ( .I1(_i_CLEFIA128_keyK _58), .I2(n14678), .O(n14679) );
  ND2HHD U9820 ( .I1(n10916), .I2(n10914), .O(n8259) );
  ND2DHD U9821 ( .I1(n10916), .I2(n10915), .O(n10917) );
  ND2CHD U9822 ( .I1(n14011), .I2(_i_CLEFIA128_rndcnt_reg _0), .O(n10500) );
  INVCHD U9823 ( .I(DOUT_62), .O(n15494) );
  INVDHD U9824 ( .I(_i_CLEFIA128_keyL _79), .O(n15186) );
  XNR2CHD U9825 ( .I1(DIN_31), .I2(_i_CLEFIA128_keyK _95), .O(n13797) );
  INVDHD U9826 ( .I(_i_CLEFIA128_keyL _15), .O(n15208) );
  INVDHD U9827 ( .I(_i_CLEFIA128_keyL _78), .O(n15409) );
  INVDHD U9828 ( .I(_i_CLEFIA128_keyL _85), .O(n15296) );
  INVCHD U9829 ( .I(DOUT_97), .O(n15271) );
  INVDHD U9830 ( .I(_i_CLEFIA128_keyL _86), .O(n15185) );
  XNR2CHD U9831 ( .I1(DIN_30), .I2(_i_CLEFIA128_keyK _94), .O(n13918) );
  INVCHD U9832 ( .I(DOUT_112), .O(n15369) );
  XOR2CHD U9833 ( .I1(DIN_31), .I2(_i_CLEFIA128_keyK _31), .O(n13794) );
  INVDHD U9834 ( .I(_i_CLEFIA128_keyL _93), .O(n15172) );
  INVDHD U9835 ( .I(_i_CLEFIA128_keyL _71), .O(n15426) );
  INVDHD U9836 ( .I(_i_CLEFIA128_keyL _92), .O(n15399) );
  INVDHD U9837 ( .I(_i_CLEFIA128_rndcnt_reg _4), .O(n7220) );
  INVDHD U9838 ( .I(_i_CLEFIA128_keyL _46), .O(n7143) );
  INVLHD U9839 ( .I(_i_CLEFIA128_keyL _36), .O(n15182) );
  INVDHD U9840 ( .I(_i_CLEFIA128_keyL _7), .O(n15398) );
  XNR2CHD U9841 ( .I1(DIN_27), .I2(_i_CLEFIA128_keyK _91), .O(n14150) );
  INVCHD U9842 ( .I(_i_CLEFIA128_keyL _106), .O(n15403) );
  INVCHD U9843 ( .I(_i_CLEFIA128_keyL _14), .O(n15407) );
  INVDHD U9844 ( .I(_i_CLEFIA128_keyL _65), .O(n15194) );
  XNR2CHD U9845 ( .I1(_i_CLEFIA128_CON_T_x _6), .I2(DOUT_102), .O(n12024) );
  INVCHD U9846 ( .I(DOUT_48), .O(n15373) );
  XOR2CHD U9847 ( .I1(DIN_27), .I2(_i_CLEFIA128_keyK _27), .O(n14147) );
  XOR2CHD U9848 ( .I1(DIN_30), .I2(_i_CLEFIA128_keyK _30), .O(n13915) );
  INVCHD U9849 ( .I(DOUT_50), .O(n14904) );
  XOR2CHD U9850 ( .I1(DIN_75), .I2(_i_CLEFIA128_keyK _43), .O(n14391) );
  INVCHD U9851 ( .I(_i_CLEFIA128_keyK _103), .O(n15469) );
  INVCHD U9852 ( .I(DOUT_43), .O(n15316) );
  INVCHD U9853 ( .I(_i_CLEFIA128_CON_T_x _8), .O(n14732) );
  XOR2CHD U9854 ( .I1(DIN_71), .I2(_i_CLEFIA128_keyK _39), .O(n15471) );
  INVCHD U9855 ( .I(DOUT_37), .O(n15043) );
  XOR2CHD U9856 ( .I1(DIN_29), .I2(_i_CLEFIA128_keyK _29), .O(n15155) );
  XOR2HHD U9857 ( .I1(_i_CLEFIA128_CON_T_x _12), .I2(DOUT_108), .O(n11864));
  XNR2CHD U9858 ( .I1(DIN_71), .I2(_i_CLEFIA128_keyK _103), .O(n15474) );
  INVCHD U9859 ( .I(_i_CLEFIA128_keyK _43), .O(n14388) );
  INVCHD U9860 ( .I(DOUT_33), .O(n15258) );
  INVDHD U9861 ( .I(_i_CLEFIA128_keyL _82), .O(n14919) );
  INVDHD U9862 ( .I(DOUT_52), .O(n14384) );
  XOR2CHD U9863 ( .I1(DIN_7), .I2(_i_CLEFIA128_keyK _7), .O(n14775) );
  INVCHD U9864 ( .I(_i_CLEFIA128_keyL _91), .O(n15128) );
  INVCHD U9865 ( .I(_i_CLEFIA128_CON_T_x _9), .O(n14736) );
  XNR2CHD U9866 ( .I1(DIN_29), .I2(_i_CLEFIA128_keyK _93), .O(n15158) );
  INVCHD U9867 ( .I(_i_CLEFIA128_keyL _75), .O(n14930) );
  XNR2CHD U9868 ( .I1(DIN_7), .I2(_i_CLEFIA128_keyK _71), .O(n14778) );
  INVCHD U9869 ( .I(DOUT_35), .O(n15055) );
  INVCHD U9870 ( .I(_i_CLEFIA128_keyL _89), .O(n14918) );
  INVCHD U9871 ( .I(DOUT_103), .O(n15483) );
  INVCHD U9872 ( .I(DOUT_41), .O(n15115) );
  INVDHD U9873 ( .I(_i_CLEFIA128_keyL _88), .O(n14972) );
  INVCHD U9874 ( .I(_i_CLEFIA128_keyK _71), .O(n14773) );
  INVCHD U9875 ( .I(_i_CLEFIA128_CON_T_x _10), .O(n14727) );
  INVCHD U9876 ( .I(DOUT_39), .O(n15475) );
  ND2CHD U9877 ( .I1(BSY), .I2(_i_CLEFIA128_keyK _122), .O(n14684) );
  XNR2CHD U9878 ( .I1(DIN_0), .I2(_i_CLEFIA128_keyK _64), .O(n15510) );
  XOR2CHD U9879 ( .I1(DIN_0), .I2(_i_CLEFIA128_keyK _0), .O(n15507) );
  INVCHD U9880 ( .I(_i_CLEFIA128_CON_T_xi _9), .O(n14731) );
  XNR2CHD U9881 ( .I1(DIN_24), .I2(_i_CLEFIA128_keyK _88), .O(n13708) );
  INVCHD U9882 ( .I(DOUT_99), .O(n15400) );
  INVCHD U9883 ( .I(_i_CLEFIA128_keyK _104), .O(n14116) );
  XOR2CHD U9884 ( .I1(DIN_24), .I2(_i_CLEFIA128_keyK _24), .O(n13705) );
  INVCHD U9885 ( .I(_i_CLEFIA128_keyK _40), .O(n14115) );
  INVCHD U9886 ( .I(_i_CLEFIA128_keyK _64), .O(n15505) );
  INVCHD U9887 ( .I(DOUT_57), .O(n15461) );
  XOR2CHD U9888 ( .I1(DIN_72), .I2(_i_CLEFIA128_keyK _40), .O(n14118) );
  INVCHD U9889 ( .I(_i_CLEFIA128_keyL _95), .O(n14979) );
  INVCHD U9890 ( .I(DOUT_106), .O(n15393) );
  INVCHD U9891 ( .I(_i_CLEFIA128_keyL _103), .O(n14957) );
  XNR2CHD U9892 ( .I1(DIN_72), .I2(_i_CLEFIA128_keyK _104), .O(n14121) );
  INVCHD U9893 ( .I(DOUT_104), .O(n15386) );
  INVDHD U9894 ( .I(_i_CLEFIA128_keyL _70), .O(n15096) );
  INVCHD U9895 ( .I(DOUT_116), .O(n14383) );
  INVCHD U9896 ( .I(_i_CLEFIA128_keyL _77), .O(n15092) );
  INVCHD U9897 ( .I(_i_CLEFIA128_CON_T_x _12), .O(n14459) );
  INVCHD U9898 ( .I(DOUT_127), .O(n15417) );
  INVCHD U9899 ( .I(DOUT_121), .O(n15462) );
  INVCHD U9900 ( .I(_i_CLEFIA128_keyK _88), .O(n13700) );
  INVCHD U9901 ( .I(DOUT_40), .O(n15385) );
  INVCHD U9902 ( .I(_i_CLEFIA128_CON_T_xi _13), .O(n14469) );
  INVCHD U9903 ( .I(DOUT_100), .O(n14814) );
  INVCHD U9904 ( .I(DOUT_102), .O(n15428) );
  XNR2CHD U9905 ( .I1(DIN_68), .I2(_i_CLEFIA128_keyK _100), .O(n13260) );
  XOR2CHD U9906 ( .I1(DIN_68), .I2(_i_CLEFIA128_keyK _36), .O(n13257) );
  INVCHD U9907 ( .I(_i_CLEFIA128_keyK _24), .O(n13699) );
  INVCHD U9908 ( .I(DOUT_114), .O(n15130) );
  INVCHD U9909 ( .I(_i_CLEFIA128_CON_T_x _0), .O(n14443) );
  INVCHD U9910 ( .I(DOUT_126), .O(n15498) );
  INVCHD U9911 ( .I(_i_CLEFIA128_keyL _124), .O(n14923) );
  INVCHD U9912 ( .I(_i_CLEFIA128_keyK _36), .O(n13255) );
  INVCHD U9913 ( .I(_i_CLEFIA128_CON_T_x _14), .O(n14449) );
  INVCHD U9914 ( .I(_i_CLEFIA128_keyK _100), .O(n13256) );
  XNR2CHD U9915 ( .I1(DIN_80), .I2(_i_CLEFIA128_keyK _112), .O(n13944) );
  INVCHD U9916 ( .I(_i_CLEFIA128_keyL _120), .O(n15415) );
  XOR2CHD U9917 ( .I1(DIN_80), .I2(_i_CLEFIA128_keyK _48), .O(n13941) );
  INVCHD U9918 ( .I(DOUT_90), .O(n9537) );
  XOR2CHD U9919 ( .I1(DIN_2), .I2(_i_CLEFIA128_keyK _2), .O(n13929) );
  INVDHD U9920 ( .I(DOUT_63), .O(n14866) );
  INVCHD U9921 ( .I(DOUT_61), .O(n15159) );
  XNR2CHD U9922 ( .I1(DIN_2), .I2(_i_CLEFIA128_keyK _66), .O(n13932) );
  INVDHD U9923 ( .I(DOUT_98), .O(n15329) );
  INVCHD U9924 ( .I(DOUT_58), .O(n14959) );
  INVCHD U9925 ( .I(DOUT_27), .O(n14139) );
  INVCHD U9926 ( .I(DOUT_59), .O(n15075) );
  INVCHD U9927 ( .I(_i_CLEFIA128_keyK _2), .O(n13922) );
  INVCHD U9928 ( .I(DOUT_60), .O(n14924) );
  INVCHD U9929 ( .I(DOUT_122), .O(n15337) );
  INVCHD U9930 ( .I(_i_CLEFIA128_keyL _105), .O(n15236) );
  INVCHD U9931 ( .I(DOUT_44), .O(n15015) );
  INVCHD U9932 ( .I(_i_CLEFIA128_keyK _27), .O(n14135) );
  INVDHD U9933 ( .I(DOUT_34), .O(n15330) );
  INVCHD U9934 ( .I(DOUT_55), .O(n15432) );
  INVCHD U9935 ( .I(_i_CLEFIA128_keyK _91), .O(n14136) );
  INVCHD U9936 ( .I(DOUT_47), .O(n15361) );
  INVCHD U9937 ( .I(DOUT_101), .O(n15030) );
  INVCHD U9938 ( .I(DOUT_54), .O(n15286) );
  INVCHD U9939 ( .I(_i_CLEFIA128_CON_T_x _2), .O(n14747) );
  INVCHD U9940 ( .I(DOUT_46), .O(n15446) );
  ND2HHD U9941 ( .I1(n8039), .I2(_i_CLEFIA128_keyK _35), .O(n9883) );
  INVCHD U9942 ( .I(_i_CLEFIA128_keyK _95), .O(n13791) );
  INVCHD U9943 ( .I(DOUT_53), .O(n14828) );
  INVCHD U9944 ( .I(_i_CLEFIA128_keyK _94), .O(n13910) );
  INVCHD U9945 ( .I(DOUT_110), .O(n15452) );
  INVCHD U9946 ( .I(DOUT_77), .O(n9592) );
  INVCHD U9947 ( .I(_i_CLEFIA128_CON_T_x _3), .O(n14753) );
  INVCHD U9948 ( .I(DOUT_45), .O(n15223) );
  INVCHD U9949 ( .I(DOUT_119), .O(n15437) );
  ND2DHD U9950 ( .I1(_i_CLEFIA128_keyL _42), .I2(_i_CLEFIA128_keyK _42), .O(n8680) );
  INVCHD U9951 ( .I(DOUT_38), .O(n15442) );
  INVCHD U9952 ( .I(DOUT_111), .O(n15360) );
  INVCHD U9953 ( .I(DOUT_36), .O(n14983) );
  INVCHD U9954 ( .I(DOUT_117), .O(n14302) );
  INVCHD U9955 ( .I(DOUT_51), .O(n15491) );
  INVCHD U9956 ( .I(_i_CLEFIA128_CON_T_reg_4 ), .O(n14739) );
  INVCHD U9957 ( .I(_i_CLEFIA128_keyK _29), .O(n15153) );
  XNR2CHD U9958 ( .I1(DIN_90), .I2(_i_CLEFIA128_keyK _122), .O(n14700) );
  INVCHD U9959 ( .I(_i_CLEFIA128_keyK _48), .O(n13936) );
  INVDHD U9960 ( .I(DOUT_49), .O(n15141) );
  XOR2CHD U9961 ( .I1(DIN_90), .I2(_i_CLEFIA128_keyK _58), .O(n14697) );
  INVCHD U9962 ( .I(_i_CLEFIA128_keyK _112), .O(n13937) );
  INVCHD U9963 ( .I(DOUT_124), .O(n14321) );
  INVCHD U9964 ( .I(DOUT_107), .O(n15317) );
  INVCHD U9965 ( .I(DOUT_108), .O(n15345) );
  INVCHD U9966 ( .I(DOUT_125), .O(n15160) );
  INVCHD U9967 ( .I(_i_CLEFIA128_CON_T_x _6), .O(n14454) );
  ND2CHD U9968 ( .I1(BSY), .I2(_i_CLEFIA128_keyK _58), .O(n14686) );
  INVCHD U9969 ( .I(DOUT_115), .O(n15488) );
  INVCHD U9970 ( .I(DOUT_109), .O(n15224) );
  INVDHD U9971 ( .I(_i_CLEFIA128_keyL _74), .O(n15301) );
  INVCHD U9972 ( .I(DOUT_42), .O(n14802) );
  XNR2CHD U9973 ( .I1(DIN_75), .I2(_i_CLEFIA128_keyK _107), .O(n14394) );
  INVCHD U9974 ( .I(DOUT_123), .O(n14291) );
  INVCHD U9975 ( .I(_i_CLEFIA128_keyK _25), .O(n15455) );
  INVCHD U9976 ( .I(_i_CLEFIA128_keyK _109), .O(n14202) );
  XNR2CHD U9977 ( .I1(DIN_3), .I2(_i_CLEFIA128_keyK _67), .O(n13272) );
  XOR2CHD U9978 ( .I1(DIN_11), .I2(_i_CLEFIA128_keyK _11), .O(n15312) );
  INVCHD U9979 ( .I(_i_CLEFIA128_keyK _45), .O(n14201) );
  INVLHD U9980 ( .I(_i_CLEFIA128_keyL _21), .O(n15137) );
  XOR2CHD U9981 ( .I1(DIN_19), .I2(_i_CLEFIA128_keyK _19), .O(n12818) );
  INVCHD U9982 ( .I(_i_CLEFIA128_keyK _111), .O(n15354) );
  XNR2CHD U9983 ( .I1(DIN_19), .I2(_i_CLEFIA128_keyK _83), .O(n12821) );
  XOR2CHD U9984 ( .I1(DIN_77), .I2(_i_CLEFIA128_keyK _45), .O(n14204) );
  XNR2CHD U9985 ( .I1(DIN_77), .I2(_i_CLEFIA128_keyK _109), .O(n14207) );
  INVCHD U9986 ( .I(_i_CLEFIA128_keyK _81), .O(n13729) );
  INVCHD U9987 ( .I(_i_CLEFIA128_keyK _17), .O(n13728) );
  XOR2CHD U9988 ( .I1(DIN_25), .I2(_i_CLEFIA128_keyK _25), .O(n15457) );
  INVCHD U9989 ( .I(_i_CLEFIA128_keyK _97), .O(n14226) );
  XNR2CHD U9990 ( .I1(DIN_25), .I2(_i_CLEFIA128_keyK _89), .O(n15460) );
  INVCHD U9991 ( .I(_i_CLEFIA128_keyK _33), .O(n14225) );
  XOR2CHD U9992 ( .I1(DIN_17), .I2(_i_CLEFIA128_keyK _17), .O(n13734) );
  INVCHD U9993 ( .I(_i_CLEFIA128_keyK _74), .O(n13971) );
  INVCHD U9994 ( .I(_i_CLEFIA128_keyK _10), .O(n13970) );
  XOR2CHD U9995 ( .I1(DIN_65), .I2(_i_CLEFIA128_keyK _33), .O(n14233) );
  XNR2CHD U9996 ( .I1(DIN_85), .I2(_i_CLEFIA128_keyK _117), .O(n14301) );
  XNR2CHD U9997 ( .I1(DIN_65), .I2(_i_CLEFIA128_keyK _97), .O(n14236) );
  XNR2CHD U9998 ( .I1(DIN_17), .I2(_i_CLEFIA128_keyK _81), .O(n13737) );
  INVCHD U9999 ( .I(_i_CLEFIA128_keyK _118), .O(n13996) );
  INVCHD U10000 ( .I(_i_CLEFIA128_keyK _102), .O(n13803) );
  INVCHD U10001 ( .I(_i_CLEFIA128_keyK _11), .O(n15309) );
  XOR2CHD U10002 ( .I1(DIN_10), .I2(_i_CLEFIA128_keyK _10), .O(n13976) );
  XOR2CHD U10003 ( .I1(DIN_12), .I2(_i_CLEFIA128_keyK _12), .O(n12888) );
  XNR2CHD U10004 ( .I1(DIN_12), .I2(_i_CLEFIA128_keyK _76), .O(n12891) );
  XNR2CHD U10005 ( .I1(DIN_10), .I2(_i_CLEFIA128_keyK _74), .O(n13979) );
  XOR2CHD U10006 ( .I1(DIN_85), .I2(_i_CLEFIA128_keyK _53), .O(n14298) );
  INVCHD U10007 ( .I(_i_CLEFIA128_keyK _75), .O(n15310) );
  XOR2CHD U10008 ( .I1(DIN_86), .I2(_i_CLEFIA128_keyK _54), .O(n13997) );
  XNR2CHD U10009 ( .I1(DIN_86), .I2(_i_CLEFIA128_keyK _118), .O(n14000) );
  XOR2CHD U10010 ( .I1(DIN_84), .I2(_i_CLEFIA128_keyK _52), .O(n14379) );
  INVCHD U10011 ( .I(_i_CLEFIA128_keyK _76), .O(n12827) );
  XNR2CHD U10012 ( .I1(DIN_84), .I2(_i_CLEFIA128_keyK _116), .O(n14382) );
  INVCHD U10013 ( .I(_i_CLEFIA128_keyK _12), .O(n12826) );
  INVCHD U10014 ( .I(_i_CLEFIA128_keyK _105), .O(n15001) );
  XOR2CHD U10015 ( .I1(DIN_87), .I2(_i_CLEFIA128_keyK _55), .O(n13770) );
  INVCHD U10016 ( .I(_i_CLEFIA128_keyK _13), .O(n15216) );
  INVCHD U10017 ( .I(_i_CLEFIA128_keyK _77), .O(n15217) );
  INVCHD U10018 ( .I(_i_CLEFIA128_keyK _21), .O(n14256) );
  XNR2CHD U10019 ( .I1(DIN_18), .I2(_i_CLEFIA128_keyK _82), .O(n13904) );
  INVCHD U10020 ( .I(_i_CLEFIA128_keyK _85), .O(n14257) );
  INVCHD U10021 ( .I(_i_CLEFIA128_keyK _53), .O(n14295) );
  INVCHD U10022 ( .I(_i_CLEFIA128_keyK _41), .O(n15000) );
  XOR2CHD U10023 ( .I1(DIN_73), .I2(_i_CLEFIA128_keyK _41), .O(n15003) );
  INVCHD U10024 ( .I(_i_CLEFIA128_keyK _117), .O(n14296) );
  XNR2CHD U10025 ( .I1(DIN_73), .I2(_i_CLEFIA128_keyK _105), .O(n15006) );
  XOR2CHD U10026 ( .I1(DIN_93), .I2(_i_CLEFIA128_keyK _61), .O(n14186) );
  XNR2CHD U10027 ( .I1(DIN_93), .I2(_i_CLEFIA128_keyK _125), .O(n14189) );
  XNR2CHD U10028 ( .I1(DIN_87), .I2(_i_CLEFIA128_keyK _119), .O(n13773) );
  INVCHD U10029 ( .I(_i_CLEFIA128_keyK _52), .O(n14376) );
  XOR2CHD U10030 ( .I1(DIN_18), .I2(_i_CLEFIA128_keyK _18), .O(n13901) );
  INVCHD U10031 ( .I(_i_CLEFIA128_keyK _125), .O(n14183) );
  XNR2CHD U10032 ( .I1(DIN_21), .I2(_i_CLEFIA128_keyK _85), .O(n14262) );
  INVCHD U10033 ( .I(_i_CLEFIA128_keyK _60), .O(n14274) );
  XOR2CHD U10034 ( .I1(DIN_21), .I2(_i_CLEFIA128_keyK _21), .O(n14259) );
  INVCHD U10035 ( .I(_i_CLEFIA128_keyK _61), .O(n14182) );
  XNR2CHD U10036 ( .I1(DIN_14), .I2(_i_CLEFIA128_keyK _78), .O(n13957) );
  INVCHD U10037 ( .I(_i_CLEFIA128_keyK _37), .O(n14211) );
  INVCHD U10038 ( .I(_i_CLEFIA128_keyK _124), .O(n14275) );
  XOR2CHD U10039 ( .I1(DIN_83), .I2(_i_CLEFIA128_keyK _51), .O(n14369) );
  XOR2CHD U10040 ( .I1(DIN_14), .I2(_i_CLEFIA128_keyK _14), .O(n13954) );
  XOR2CHD U10041 ( .I1(DIN_81), .I2(_i_CLEFIA128_keyK _49), .O(n14158) );
  XNR2CHD U10042 ( .I1(DIN_83), .I2(_i_CLEFIA128_keyK _115), .O(n14372) );
  XNR2CHD U10043 ( .I1(DIN_81), .I2(_i_CLEFIA128_keyK _113), .O(n14161) );
  INVCHD U10044 ( .I(_i_CLEFIA128_keyK _78), .O(n13950) );
  XOR2CHD U10045 ( .I1(DIN_67), .I2(_i_CLEFIA128_keyK _35), .O(n14334) );
  INVCHD U10046 ( .I(_i_CLEFIA128_keyK _5), .O(n14241) );
  XNR2CHD U10047 ( .I1(DIN_6), .I2(_i_CLEFIA128_keyK _70), .O(n14022) );
  INVCHD U10048 ( .I(_i_CLEFIA128_keyK _35), .O(n14325) );
  INVCHD U10049 ( .I(DOUT_105), .O(n15106) );
  INVCHD U10050 ( .I(_i_CLEFIA128_keyK _70), .O(n14012) );
  INVCHD U10051 ( .I(_i_CLEFIA128_keyL _112), .O(n15249) );
  INVCHD U10052 ( .I(_i_CLEFIA128_keyK _120), .O(n14041) );
  INVCHD U10053 ( .I(_i_CLEFIA128_keyK _56), .O(n14040) );
  XNR2CHD U10054 ( .I1(DIN_8), .I2(_i_CLEFIA128_keyK _72), .O(n15384) );
  INVCHD U10055 ( .I(_i_CLEFIA128_keyK _68), .O(n10304) );
  INVCHD U10056 ( .I(_i_CLEFIA128_keyK _4), .O(n10303) );
  XOR2CHD U10057 ( .I1(DIN_5), .I2(_i_CLEFIA128_keyK _5), .O(n14249) );
  XOR2CHD U10058 ( .I1(DIN_8), .I2(_i_CLEFIA128_keyK _8), .O(n15381) );
  XNR2CHD U10059 ( .I1(DIN_5), .I2(_i_CLEFIA128_keyK _69), .O(n14252) );
  XOR2CHD U10060 ( .I1(DIN_88), .I2(_i_CLEFIA128_keyK _56), .O(n14094) );
  INVCHD U10061 ( .I(_i_CLEFIA128_keyK _8), .O(n15378) );
  INVCHD U10062 ( .I(_i_CLEFIA128_keyK _72), .O(n15379) );
  INVCHD U10063 ( .I(_i_CLEFIA128_keyK _110), .O(n14027) );
  XNR2CHD U10064 ( .I1(DIN_9), .I2(_i_CLEFIA128_keyK _73), .O(n13760) );
  INVCHD U10065 ( .I(_i_CLEFIA128_keyK _101), .O(n14212) );
  XNR2CHD U10066 ( .I1(DIN_88), .I2(_i_CLEFIA128_keyK _120), .O(n14097) );
  XOR2CHD U10067 ( .I1(DIN_9), .I2(_i_CLEFIA128_keyK _9), .O(n13757) );
  XNR2CHD U10068 ( .I1(DIN_13), .I2(_i_CLEFIA128_keyK _77), .O(n15222) );
  INVCHD U10069 ( .I(_i_CLEFIA128_keyK _1), .O(n13713) );
  XOR2CHD U10070 ( .I1(DIN_13), .I2(_i_CLEFIA128_keyK _13), .O(n15219) );
  INVCHD U10071 ( .I(_i_CLEFIA128_keyK _9), .O(n13752) );
  XOR2CHD U10072 ( .I1(DIN_6), .I2(_i_CLEFIA128_keyK _6), .O(n14019) );
  INVCHD U10073 ( .I(_i_CLEFIA128_keyK _73), .O(n9974) );
  XNR2CHD U10074 ( .I1(DIN_16), .I2(_i_CLEFIA128_keyK _80), .O(n13785) );
  XOR2CHD U10075 ( .I1(DIN_16), .I2(_i_CLEFIA128_keyK _16), .O(n13782) );
  XOR2CHD U10076 ( .I1(DIN_1), .I2(_i_CLEFIA128_keyK _1), .O(n13720) );
  XNR2CHD U10077 ( .I1(DIN_1), .I2(_i_CLEFIA128_keyK _65), .O(n13723) );
  INVCHD U10078 ( .I(_i_CLEFIA128_keyK _50), .O(n13041) );
  INVCHD U10079 ( .I(_i_CLEFIA128_keyK _119), .O(n13766) );
  INVCHD U10080 ( .I(_i_CLEFIA128_keyK _16), .O(n13777) );
  INVLHD U10081 ( .I(_i_CLEFIA128_keyL _1), .O(n15209) );
  INVCHD U10082 ( .I(_i_CLEFIA128_keyK _34), .O(n15322) );
  INVCHD U10083 ( .I(_i_CLEFIA128_keyK _98), .O(n15323) );
  XNR2CHD U10084 ( .I1(DIN_66), .I2(_i_CLEFIA128_keyK _98), .O(n15328) );
  XOR2CHD U10085 ( .I1(DIN_66), .I2(_i_CLEFIA128_keyK _34), .O(n15325) );
  XOR2CHD U10086 ( .I1(DIN_4), .I2(_i_CLEFIA128_keyK _4), .O(n10918) );
  XOR2CHD U10087 ( .I1(DIN_20), .I2(_i_CLEFIA128_keyK _20), .O(n10929) );
  XNR2CHD U10088 ( .I1(DIN_4), .I2(_i_CLEFIA128_keyK _68), .O(n10921) );
  XNR2CHD U10089 ( .I1(DIN_20), .I2(_i_CLEFIA128_keyK _84), .O(n10932) );
  XNR2CHD U10090 ( .I1(DIN_79), .I2(_i_CLEFIA128_keyK _111), .O(n15359) );
  XNR2CHD U10091 ( .I1(DIN_69), .I2(_i_CLEFIA128_keyK _101), .O(n14221) );
  XOR2CHD U10092 ( .I1(DIN_69), .I2(_i_CLEFIA128_keyK _37), .O(n14218) );
  INVCHD U10093 ( .I(_i_CLEFIA128_keyK _20), .O(n10935) );
  INVCHD U10094 ( .I(_i_CLEFIA128_keyK _83), .O(n12595) );
  INVCHD U10095 ( .I(_i_CLEFIA128_keyK _19), .O(n12594) );
  XOR2CHD U10096 ( .I1(DIN_82), .I2(_i_CLEFIA128_keyK _50), .O(n13042) );
  XNR2CHD U10097 ( .I1(DIN_82), .I2(_i_CLEFIA128_keyK _114), .O(n13045) );
  XOR2CHD U10098 ( .I1(DIN_79), .I2(_i_CLEFIA128_keyK _47), .O(n15356) );
  XNR2CHD U10099 ( .I1(DIN_78), .I2(_i_CLEFIA128_keyK _110), .O(n14036) );
  XNR2CHD U10100 ( .I1(DIN_11), .I2(_i_CLEFIA128_keyK _75), .O(n15315) );
  XOR2CHD U10101 ( .I1(DIN_3), .I2(_i_CLEFIA128_keyK _3), .O(n13269) );
  XOR2CHD U10102 ( .I1(DIN_78), .I2(_i_CLEFIA128_keyK _46), .O(n14033) );
  INVCHD U10103 ( .I(_i_CLEFIA128_keyK _87), .O(n13882) );
  INVCHD U10104 ( .I(_i_CLEFIA128_keyK _127), .O(n14755) );
  XOR2CHD U10105 ( .I1(DIN_26), .I2(_i_CLEFIA128_keyK _26), .O(n13873) );
  INVCHD U10106 ( .I(_i_CLEFIA128_keyK _26), .O(n13869) );
  INVCHD U10107 ( .I(_i_CLEFIA128_keyK _90), .O(n13870) );
  INVCHD U10108 ( .I(DOUT_32), .O(n15511) );
  XNR2CHD U10109 ( .I1(DIN_91), .I2(_i_CLEFIA128_keyK _123), .O(n14290) );
  XOR2CHD U10110 ( .I1(DIN_91), .I2(_i_CLEFIA128_keyK _59), .O(n14287) );
  INVCHD U10111 ( .I(_i_CLEFIA128_keyK _18), .O(n13893) );
  XOR2CHD U10112 ( .I1(DIN_23), .I2(_i_CLEFIA128_keyK _23), .O(n13886) );
  INVCHD U10113 ( .I(_i_CLEFIA128_keyK _82), .O(n13894) );
  XNR2CHD U10114 ( .I1(DIN_76), .I2(_i_CLEFIA128_keyK _108), .O(n14311) );
  INVCHD U10115 ( .I(_i_CLEFIA128_keyK _57), .O(n14885) );
  XOR2CHD U10116 ( .I1(DIN_89), .I2(_i_CLEFIA128_keyK _57), .O(n14887) );
  XNR2CHD U10117 ( .I1(DIN_23), .I2(_i_CLEFIA128_keyK _87), .O(n13889) );
  INVCHD U10118 ( .I(_i_CLEFIA128_keyL _104), .O(n15274) );
  XNR2CHD U10119 ( .I1(DIN_64), .I2(_i_CLEFIA128_keyK _96), .O(n14131) );
  INVCHD U10120 ( .I(_i_CLEFIA128_keyK _79), .O(n14785) );
  XOR2CHD U10121 ( .I1(DIN_76), .I2(_i_CLEFIA128_keyK _44), .O(n14308) );
  INVCHD U10122 ( .I(_i_CLEFIA128_keyK _49), .O(n14154) );
  XNR2CHD U10123 ( .I1(DIN_26), .I2(_i_CLEFIA128_keyK _90), .O(n13876) );
  XOR2CHD U10124 ( .I1(DIN_95), .I2(_i_CLEFIA128_keyK _63), .O(n14757) );
  INVCHD U10125 ( .I(_i_CLEFIA128_keyL _90), .O(n15270) );
  XOR2CHD U10126 ( .I1(DIN_64), .I2(_i_CLEFIA128_keyK _32), .O(n14128) );
  INVCHD U10127 ( .I(_i_CLEFIA128_keyK _113), .O(n14155) );
  XNR2CHD U10128 ( .I1(DIN_74), .I2(_i_CLEFIA128_keyK _106), .O(n14357) );
  XOR2CHD U10129 ( .I1(DIN_15), .I2(_i_CLEFIA128_keyK _15), .O(n14787) );
  INVCHD U10130 ( .I(DOUT_96), .O(n15514) );
  XOR2CHD U10131 ( .I1(DIN_74), .I2(_i_CLEFIA128_keyK _42), .O(n14354) );
  XNR2CHD U10132 ( .I1(DIN_15), .I2(_i_CLEFIA128_keyK _79), .O(n14790) );
  XNR2CHD U10133 ( .I1(DIN_94), .I2(_i_CLEFIA128_keyK _126), .O(n13695) );
  XNR2CHD U10134 ( .I1(DIN_28), .I2(_i_CLEFIA128_keyK _92), .O(n14320) );
  INVCHD U10135 ( .I(_i_CLEFIA128_keyL _83), .O(n15293) );
  XNR2CHD U10136 ( .I1(DIN_89), .I2(_i_CLEFIA128_keyK _121), .O(n14890) );
  INVCHD U10137 ( .I(_i_CLEFIA128_keyK _42), .O(n14349) );
  INVCHD U10138 ( .I(_i_CLEFIA128_keyK _32), .O(n14125) );
  XNR2CHD U10139 ( .I1(DIN_95), .I2(_i_CLEFIA128_keyK _127), .O(n14760) );
  INVCHD U10140 ( .I(_i_CLEFIA128_keyK _44), .O(n14306) );
  XOR2CHD U10141 ( .I1(DIN_28), .I2(_i_CLEFIA128_keyK _28), .O(n14317) );
  INVCHD U10142 ( .I(_i_CLEFIA128_keyK _86), .O(n13985) );
  INVCHD U10143 ( .I(_i_CLEFIA128_keyK _96), .O(n14126) );
  INVDHD U10144 ( .I(_i_CLEFIA128_keyL _66), .O(n15344) );
  INVDHD U10145 ( .I(_i_CLEFIA128_keyL _76), .O(n15061) );
  INVDHD U10146 ( .I(_i_CLEFIA128_keyL _30), .O(n15046) );
  INVCHD U10147 ( .I(_i_CLEFIA128_keyK _123), .O(n14285) );
  XNR2CHD U10148 ( .I1(DIN_92), .I2(_i_CLEFIA128_keyK _124), .O(n14280) );
  INVDHD U10149 ( .I(_i_CLEFIA128_keyL _94), .O(n15050) );
  INVCHD U10150 ( .I(_i_CLEFIA128_keyK _106), .O(n14350) );
  XNR2CHD U10151 ( .I1(DIN_70), .I2(_i_CLEFIA128_keyK _102), .O(n13857) );
  XOR2CHD U10152 ( .I1(DIN_94), .I2(_i_CLEFIA128_keyK _62), .O(n13692) );
  XNR2CHD U10153 ( .I1(_i_CLEFIA128_CON_T_x _8), .I2(DOUT_47), .O(n8405) );
  INVCHD U10154 ( .I(_i_CLEFIA128_keyK _92), .O(n14316) );
  INVCHD U10155 ( .I(_i_CLEFIA128_keyK _126), .O(n13571) );
  XOR2CHD U10156 ( .I1(DIN_92), .I2(_i_CLEFIA128_keyK _60), .O(n14277) );
  XOR2CHD U10157 ( .I1(DIN_22), .I2(_i_CLEFIA128_keyK _22), .O(n13988) );
  INVCHD U10158 ( .I(_i_CLEFIA128_keyK _115), .O(n14362) );
  XNR2CHD U10159 ( .I1(DIN_22), .I2(_i_CLEFIA128_keyK _86), .O(n13991) );
  INVDHD U10160 ( .I(_i_CLEFIA128_keyL _87), .O(n15036) );
  INVCHD U10161 ( .I(_i_CLEFIA128_keyK _59), .O(n14284) );
  INVCHD U10162 ( .I(_i_CLEFIA128_keyK _51), .O(n14361) );
  ND2DHD U10163 ( .I1(_i_CLEFIA128_keyL _94), .I2(_i_CLEFIA128_keyK _94), .O(n7532) );
  INVCHD U10164 ( .I(_i_CLEFIA128_keyK _108), .O(n14307) );
  XOR2CHD U10165 ( .I1(DIN_70), .I2(_i_CLEFIA128_keyK _38), .O(n13854) );
  INVLHD U10166 ( .I(_i_CLEFIA128_keyL _18), .O(n14950) );
  INVCHD U10167 ( .I(DOUT_118), .O(n15251) );
  INVCHD U10168 ( .I(_i_CLEFIA128_keyK _28), .O(n14315) );
  NR2GHD U10169 ( .I1(MODE_0), .I2(n10913), .O(n10914) );
  AN2HHD U10170 ( .I1(n12416), .I2(n13458), .O(n9859) );
  NR2GHD U10171 ( .I1(n7424), .I2(n12415), .O(n9090) );
  ND2KHD U10172 ( .I1(n11274), .I2(n9087), .O(n12486) );
  ND2KHD U10173 ( .I1(n8115), .I2(n6831), .O(n7776) );
  INVNHD U10174 ( .I(n7775), .O(n11713) );
  ND2KHD U10175 ( .I1(n9185), .I2(n14083), .O(n8029) );
  NR2GHD U10176 ( .I1(n7614), .I2(n7615), .O(n7428) );
  OA12HHD U10177 ( .B1(n10056), .B2(n13816), .A1(n13817), .O(n10055) );
  ND3EHD U10178 ( .I1(n8701), .I2(n12303), .I3(n12297), .O(n13816) );
  INVQHD U10179 ( .I(_i_CLEFIA128_keyL _67), .O(n15304) );
  ND3EHD U10180 ( .I1(n7681), .I2(n8430), .I3(n8247), .O(n11361) );
  NR2GHD U10181 ( .I1(n7694), .I2(n8862), .O(n7693) );
  ND2KHD U10182 ( .I1(n9184), .I2(n8210), .O(n11852) );
  ND3EHD U10183 ( .I1(n12804), .I2(n8685), .I3(n12805), .O(n8635) );
  NR2GHD U10184 ( .I1(n7880), .I2(n7246), .O(n8685) );
  ND2KHD U10185 ( .I1(n10664), .I2(n7168), .O(n10792) );
  ND3EHD U10186 ( .I1(n12913), .I2(n10228), .I3(n10131), .O(n7046) );
  ND3EHD U10187 ( .I1(n8994), .I2(n7047), .I3(n9172), .O(n9821) );
  ND3EHD U10188 ( .I1(n12406), .I2(n12405), .I3(n13120), .O(n12407) );
  BUFIHD U10189 ( .I(n8115), .O(n7934) );
  NR2EHD U10190 ( .I1(n8648), .I2(n8649), .O(n8647) );
  ND2HHD U10191 ( .I1(n9406), .I2(n13051), .O(n7765) );
  NR2IHD U10192 ( .I1(n6907), .I2(n9946), .O(n9406) );
  ND2KHD U10193 ( .I1(n8078), .I2(n9628), .O(n13085) );
  NR2CHD U10194 ( .I1(n12059), .I2(n12404), .O(n12061) );
  NR2GHD U10195 ( .I1(n10443), .I2(n10737), .O(n9855) );
  ND2HHD U10196 ( .I1(n12847), .I2(n8511), .O(n8958) );
  ND3EHD U10197 ( .I1(n9725), .I2(n11478), .I3(n11477), .O(n11481) );
  ND3EHD U10198 ( .I1(n7196), .I2(n12590), .I3(n10064), .O(n7131) );
  ND3EHD U10199 ( .I1(n7782), .I2(n7780), .I3(n7781), .O(n7727) );
  NR2GHD U10200 ( .I1(n11476), .I2(n11475), .O(n11477) );
  OA12HHD U10201 ( .B1(n9389), .B2(n11128), .A1(n8328), .O(n9009) );
  XNR2KHD U10202 ( .I1(n10231), .I2(n10230), .O(n9389) );
  INVLHD U10203 ( .I(n10259), .O(n7132) );
  INVCKIHD U10204 ( .I(n8853), .O(n8852) );
  AN2HHD U10205 ( .I1(n13366), .I2(n12955), .O(n8433) );
  ND3EHD U10206 ( .I1(n11986), .I2(n11985), .I3(n7389), .O(n11987) );
  ND2KHD U10207 ( .I1(n12558), .I2(n11511), .O(n11406) );
  ND3EHD U10208 ( .I1(n12313), .I2(n13660), .I3(n13511), .O(n9032) );
  NR2IHD U10209 ( .I1(n8856), .I2(n7023), .O(n12313) );
  ND2HHD U10210 ( .I1(n8039), .I2(_i_CLEFIA128_keyK _106), .O(n11876) );
  ND2KHD U10211 ( .I1(n9639), .I2(n13195), .O(n7870) );
  ND2KHD U10212 ( .I1(n9580), .I2(n11995), .O(n9639) );
  ND2KHD U10213 ( .I1(n9422), .I2(n9628), .O(n9667) );
  ND2KHD U10214 ( .I1(n7254), .I2(n7386), .O(n7859) );
  ND3EHD U10215 ( .I1(n12582), .I2(n11358), .I3(n7307), .O(n7493) );
  ND2HHD U10216 ( .I1(n10250), .I2(n9894), .O(n9451) );
  INVMHD U10217 ( .I(n9110), .O(n11175) );
  XOR2HHD U10218 ( .I1(n9870), .I2(n7055), .O(n8074) );
  INVNHD U10219 ( .I(_i_CLEFIA128_keyL _9), .O(n15352) );
  ND2HHD U10220 ( .I1(n10066), .I2(n10065), .O(n9685) );
  INVGHD U10221 ( .I(n7056), .O(n12343) );
  ND3EHD U10222 ( .I1(n13401), .I2(n12431), .I3(n12361), .O(n7056) );
  ND2KHD U10223 ( .I1(n9678), .I2(n9239), .O(n13029) );
  ND2HHD U10224 ( .I1(n8463), .I2(n12725), .O(n10054) );
  OAI12CHD U10225 ( .B1(n7613), .B2(n11129), .A1(n7057), .O(n6195) );
  AN2HHD U10226 ( .I1(n8075), .I2(n14671), .O(n7057) );
  ND2KHD U10227 ( .I1(n10425), .I2(n12704), .O(n10946) );
  AN2EHD U10228 ( .I1(n7835), .I2(n13659), .O(n13677) );
  NR2IHD U10229 ( .I1(n9825), .I2(n9826), .O(n7838) );
  AN2HHD U10230 ( .I1(n13426), .I2(n13425), .O(n8266) );
  INVCKIHD U10231 ( .I(n8212), .O(n8137) );
  ND2KHD U10232 ( .I1(n7866), .I2(n10326), .O(n9329) );
  INVGHD U10233 ( .I(n7059), .O(n10592) );
  ND3EHD U10234 ( .I1(n10591), .I2(n8782), .I3(n8409), .O(n7059) );
  ND3EHD U10235 ( .I1(n12775), .I2(n12777), .I3(n12776), .O(n12779) );
  AN2HHD U10236 ( .I1(n11493), .I2(n11339), .O(n12777) );
  ND3EHD U10237 ( .I1(n11491), .I2(n11382), .I3(n8452), .O(n8015) );
  NR2IHD U10238 ( .I1(n10426), .I2(n7783), .O(n9384) );
  OR3HHD U10239 ( .I1(n11516), .I2(n11515), .I3(n11514), .O(n11517) );
  ND3EHD U10240 ( .I1(n8101), .I2(n11337), .I3(n11358), .O(n11515) );
  OR2EHD U10241 ( .I1(n15267), .I2(n11921), .O(n7060) );
  ND2HHD U10242 ( .I1(n11925), .I2(n15289), .O(n7062) );
  AN2HHD U10243 ( .I1(n8116), .I2(n11027), .O(n7097) );
  ND2DHD U10244 ( .I1(n7186), .I2(n7043), .O(n7243) );
  ND2HHD U10245 ( .I1(n7109), .I2(n12586), .O(n12587) );
  NR2IHD U10246 ( .I1(n11519), .I2(n11518), .O(n9073) );
  ND3EHD U10247 ( .I1(n8698), .I2(n9392), .I3(n8999), .O(n7064) );
  INVQHD U10248 ( .I(_i_CLEFIA128_keyK _84), .O(n9132) );
  ND2HHD U10249 ( .I1(n12681), .I2(n10888), .O(n10034) );
  NR2GHD U10250 ( .I1(n7728), .I2(n7065), .O(n8956) );
  ND2HHD U10251 ( .I1(n8233), .I2(n9459), .O(n7065) );
  ND2HHD U10252 ( .I1(n7068), .I2(n8568), .O(n14490) );
  OAI12CHD U10253 ( .B1(n10854), .B2(n8873), .A1(n10853), .O(n7068) );
  ND3EHD U10254 ( .I1(n8525), .I2(n7289), .I3(n10469), .O(n8522) );
  ND2KHD U10255 ( .I1(n7180), .I2(n8447), .O(n7312) );
  ND2KHD U10256 ( .I1(n9841), .I2(n7397), .O(n11020) );
  ND2KHD U10257 ( .I1(n12618), .I2(n11254), .O(n7138) );
  ND3EHD U10258 ( .I1(n12618), .I2(n12521), .I3(n12635), .O(n9585) );
  ND2KHD U10259 ( .I1(n10802), .I2(n9659), .O(n12618) );
  NR2CHD U10260 ( .I1(n13026), .I2(n13032), .O(n9253) );
  OR3HHD U10261 ( .I1(n12801), .I2(n12800), .I3(n12799), .O(n12802) );
  ND2KHD U10262 ( .I1(n10219), .I2(n7723), .O(n12674) );
  XNR3EHD U10263 ( .I1(n7956), .I2(n6815), .I3(n7955), .O(n9374) );
  ND2DHD U10264 ( .I1(n11910), .I2(n11909), .O(n11927) );
  ND2KHD U10265 ( .I1(n9597), .I2(n9183), .O(n8253) );
  ND2HHD U10266 ( .I1(n8797), .I2(_i_CLEFIA128_keyK _32), .O(n7069) );
  ND3EHD U10267 ( .I1(n7070), .I2(n14936), .I3(_i_CLEFIA128_rndcnt_reg _0), .O(n11584) );
  ND2HHD U10268 ( .I1(n7219), .I2(_i_CLEFIA128_keyK _60), .O(n7070) );
  ND2HHD U10269 ( .I1(n8508), .I2(n12692), .O(n8809) );
  NR2GHD U10270 ( .I1(n8447), .I2(n7180), .O(n10247) );
  ND2HHD U10271 ( .I1(n6557), .I2(n11130), .O(n8169) );
  ND2KHD U10272 ( .I1(n8204), .I2(n9183), .O(n13470) );
  OR3HHD U10273 ( .I1(n9748), .I2(n11414), .I3(n7661), .O(n12565) );
  ND2HHD U10274 ( .I1(n11119), .I2(n7146), .O(n11414) );
  ND2HHD U10275 ( .I1(n13440), .I2(n12431), .O(n7844) );
  NR2IHD U10276 ( .I1(n10431), .I2(n9444), .O(n7474) );
  NR2GHD U10277 ( .I1(n11483), .I2(n9036), .O(n9796) );
  ND2HHD U10278 ( .I1(n9599), .I2(n12506), .O(n9598) );
  XNR3EHD U10279 ( .I1(n7072), .I2(n14803), .I3(n8766), .O(n8586) );
  XOR2HHD U10280 ( .I1(n7073), .I2(n10018), .O(n7072) );
  NR2GHD U10281 ( .I1(n8811), .I2(n8810), .O(n8808) );
  ND2KHD U10282 ( .I1(n9042), .I2(n9330), .O(n7477) );
  ND3EHD U10283 ( .I1(n10579), .I2(n10580), .I3(_i_CLEFIA128_state_reg _1), .O(n10581) );
  ND2KHD U10284 ( .I1(n9830), .I2(n7872), .O(n9102) );
  AN2HHD U10285 ( .I1(n15137), .I2(_i_CLEFIA128_rndcnt_reg _0), .O(n8367) );
  ND2KHD U10286 ( .I1(n7723), .I2(n12829), .O(n9735) );
  ND2KHD U10287 ( .I1(n9184), .I2(n6837), .O(n14083) );
  NR2GHD U10288 ( .I1(n10439), .I2(n10284), .O(n10440) );
  ND3EHD U10289 ( .I1(n9703), .I2(n10438), .I3(n8337), .O(n10284) );
  ND3EHD U10290 ( .I1(n11531), .I2(n11443), .I3(n12450), .O(n9901) );
  AN2HHD U10291 ( .I1(n12486), .I2(n10624), .O(n10625) );
  ND2KHD U10292 ( .I1(n10794), .I2(n10179), .O(n8235) );
  ND3EHD U10293 ( .I1(n10225), .I2(n11840), .I3(n9568), .O(n8186) );
  NR2IHD U10294 ( .I1(n9566), .I2(n9565), .O(n8076) );
  NR2IHD U10295 ( .I1(n7075), .I2(n7074), .O(n8023) );
  INVGHD U10296 ( .I(n8024), .O(n7075) );
  NR2EHD U10297 ( .I1(n13103), .I2(n8645), .O(n8644) );
  OA12HHD U10298 ( .B1(n7910), .B2(n12201), .A1(n14049), .O(n7909) );
  NR2IHD U10299 ( .I1(n13058), .I2(n11832), .O(n7076) );
  ND2KHD U10300 ( .I1(n11614), .I2(n8800), .O(n11832) );
  BUFEHD U10301 ( .I(n7394), .O(n7078) );
  NR2GHD U10302 ( .I1(n10640), .I2(n10639), .O(n10641) );
  INVKHD U10303 ( .I(n9612), .O(n10143) );
  OAI112BHD U10304 ( .C1(n9697), .C2(n13853), .A1(n7079), .B1(n13860), .O(n6152) );
  ND2HHD U10305 ( .I1(n9697), .I2(n13852), .O(n7079) );
  OR3HHD U10306 ( .I1(n12965), .I2(n13017), .I3(n12964), .O(n12974) );
  BUFKHD U10307 ( .I(n9406), .O(n7080) );
  ND2KHD U10308 ( .I1(n10794), .I2(n10668), .O(n12651) );
  ND2KHD U10309 ( .I1(n7204), .I2(n7203), .O(n8159) );
  INVGHD U10310 ( .I(n13506), .O(n11796) );
  ND2HHD U10311 ( .I1(n7084), .I2(n7444), .O(n7443) );
  NR2EHD U10312 ( .I1(n9524), .I2(n7341), .O(n10882) );
  OAI112BHD U10313 ( .C1(n7613), .C2(n15513), .A1(n8301), .B1(n9616), .O(n6163) );
  ND3EHD U10314 ( .I1(n10454), .I2(n8020), .I3(n8019), .O(n7086) );
  XNR2KHD U10315 ( .I1(n7088), .I2(n8586), .O(n15171) );
  XOR2HHD U10316 ( .I1(n14805), .I2(n14804), .O(n7088) );
  NR2IHD U10317 ( .I1(n8507), .I2(n8505), .O(n8504) );
  ND2KHD U10318 ( .I1(n13690), .I2(n9820), .O(n9816) );
  ND2HHD U10319 ( .I1(n7091), .I2(n7090), .O(n11420) );
  INVCKIHD U10320 ( .I(n9143), .O(n7090) );
  ND2KHD U10321 ( .I1(n7093), .I2(n7092), .O(n10191) );
  INVJHD U10322 ( .I(n7044), .O(n7092) );
  ND2KHD U10323 ( .I1(n11766), .I2(n6837), .O(n13487) );
  ND2HHD U10324 ( .I1(n7095), .I2(n7094), .O(n7436) );
  NR2GHD U10325 ( .I1(n8435), .I2(n7989), .O(n7094) );
  XOR2HHD U10326 ( .I1(n14213), .I2(n7506), .O(n7505) );
  XNR2KHD U10327 ( .I1(n9543), .I2(n8898), .O(n14525) );
  INVNHD U10328 ( .I(n9644), .O(n8938) );
  INVGHD U10329 ( .I(n11661), .O(n7545) );
  AN3HHD U10330 ( .I1(n9011), .I2(n7491), .I3(n11359), .O(n7490) );
  ND2HHD U10331 ( .I1(n8824), .I2(n7434), .O(n7432) );
  ND2HHD U10332 ( .I1(n8899), .I2(n11963), .O(n8824) );
  ND2DHD U10333 ( .I1(n15307), .I2(n8283), .O(n8703) );
  XNR2KHD U10334 ( .I1(n14333), .I2(n7837), .O(n15307) );
  OA13EHD U10335 ( .B1(n13675), .B2(n13676), .B3(n13674), .A1(n8294), .O(n13689) );
  ND2HHD U10336 ( .I1(n7831), .I2(n11130), .O(n15495) );
  AN2HHD U10337 ( .I1(n7228), .I2(_i_CLEFIA128_state_reg _1), .O(n7096) );
  NR2GHD U10338 ( .I1(n7098), .I2(n7097), .O(n11028) );
  INVGHD U10339 ( .I(n7578), .O(n7536) );
  ND2HHD U10340 ( .I1(n7420), .I2(n10738), .O(n12877) );
  ND3CHD U10341 ( .I1(n8425), .I2(n12674), .I3(n12688), .O(n10815) );
  BUFQHD U10342 ( .I(n10739), .O(n10123) );
  ND3EHD U10343 ( .I1(n8951), .I2(n8950), .I3(n8949), .O(n7100) );
  AN2HHD U10344 ( .I1(n12768), .I2(n12778), .O(n12575) );
  ND2KHD U10345 ( .I1(n7313), .I2(n7314), .O(n7180) );
  NR2GHD U10346 ( .I1(n10120), .I2(n7101), .O(n10119) );
  ND3EHD U10347 ( .I1(n12449), .I2(n9237), .I3(n9128), .O(n7101) );
  BUFEHD U10348 ( .I(n7783), .O(n7102) );
  NR2IHD U10349 ( .I1(n7040), .I2(n10972), .O(n8739) );
  ND2KHD U10350 ( .I1(n9581), .I2(n7420), .O(n8194) );
  ND2HHD U10351 ( .I1(n8221), .I2(n6919), .O(n11654) );
  NR2EHD U10352 ( .I1(n10777), .I2(n7134), .O(n10780) );
  NR2IHD U10353 ( .I1(n8207), .I2(n7879), .O(n8991) );
  INVNHD U10354 ( .I(n8130), .O(n8224) );
  NR2IHD U10355 ( .I1(n9174), .I2(n9171), .O(n9169) );
  OR3HHD U10356 ( .I1(n10801), .I2(n10877), .I3(n10671), .O(n10678) );
  NR2IHD U10357 ( .I1(n9036), .I2(n11475), .O(n11348) );
  ND2KHD U10358 ( .I1(n9817), .I2(n8258), .O(n9715) );
  XNR2KHD U10359 ( .I1(n7868), .I2(n12445), .O(n14194) );
  ND2KHD U10360 ( .I1(n7198), .I2(n10266), .O(n7775) );
  XNR2KHD U10361 ( .I1(n14227), .I2(n8830), .O(n14695) );
  OA12HHD U10362 ( .B1(n9389), .B2(n11129), .A1(n8241), .O(n9077) );
  OA13HHD U10363 ( .B1(n12096), .B2(n6533), .B3(n12095), .A1(n13835), .O(n9000) );
  NR2GHD U10364 ( .I1(n7728), .I2(n10451), .O(n7730) );
  ND2HHD U10365 ( .I1(n8875), .I2(n11130), .O(n9021) );
  NR2EHD U10366 ( .I1(n9434), .I2(n8265), .O(n9740) );
  AN2HHD U10367 ( .I1(n12743), .I2(n12765), .O(n11367) );
  ND3EHD U10368 ( .I1(n7660), .I2(n11408), .I3(n7659), .O(n7658) );
  XOR2HHD U10369 ( .I1(DOUT_28), .I2(n7195), .O(n9955) );
  ND2KHD U10370 ( .I1(n9624), .I2(n9076), .O(n7195) );
  NR2IHD U10371 ( .I1(n7698), .I2(n12081), .O(n7696) );
  ND2KHD U10372 ( .I1(n12264), .I2(n9206), .O(n12000) );
  ND3EHD U10373 ( .I1(n7108), .I2(n7201), .I3(n11980), .O(n8158) );
  INVJHD U10374 ( .I(n8159), .O(n7108) );
  AN2HHD U10375 ( .I1(n10644), .I2(n9766), .O(n9575) );
  NR2IHD U10376 ( .I1(n8798), .I2(n13714), .O(n8001) );
  ND2DHD U10377 ( .I1(n10661), .I2(n7507), .O(n11225) );
  ND3EHD U10378 ( .I1(n9117), .I2(n13009), .I3(n13008), .O(n13010) );
  NR2GHD U10379 ( .I1(n11409), .I2(n12574), .O(n10052) );
  INVGHD U10380 ( .I(n7551), .O(n12258) );
  INVGHD U10381 ( .I(n11079), .O(n11074) );
  ND2HHD U10382 ( .I1(n8797), .I2(_i_CLEFIA128_keyK _90), .O(n10321) );
  ND2HHD U10383 ( .I1(n7139), .I2(n13004), .O(n13007) );
  OAI12CHD U10384 ( .B1(n8116), .B2(n8180), .A1(n9898), .O(n11091) );
  INVNHD U10385 ( .I(n8775), .O(n10973) );
  INVCKIHD U10386 ( .I(n8100), .O(n7491) );
  ND3EHD U10387 ( .I1(n8251), .I2(n11232), .I3(n7018), .O(n10368) );
  ND2DHD U10388 ( .I1(n10528), .I2(n8469), .O(n10529) );
  ND3EHD U10389 ( .I1(n10532), .I2(n10531), .I3(n10530), .O(n11125) );
  NR2GHD U10390 ( .I1(n11839), .I2(n11840), .O(n11631) );
  ND2HHD U10391 ( .I1(n12610), .I2(n7375), .O(n10807) );
  ND2KHD U10392 ( .I1(n10802), .I2(n10874), .O(n12610) );
  INVGHD U10393 ( .I(n13470), .O(n7895) );
  OAI112BHD U10394 ( .C1(n7082), .C2(n13928), .A1(n7111), .B1(n13935), .O(n6125) );
  INVGHD U10395 ( .I(n8060), .O(n13220) );
  ND2KHD U10396 ( .I1(n14427), .I2(BSY), .O(n11129) );
  ND2HHD U10397 ( .I1(n9747), .I2(n12268), .O(n12005) );
  XNR2KHD U10398 ( .I1(n14345), .I2(n8796), .O(n7231) );
  ND3EHD U10399 ( .I1(n7921), .I2(n7920), .I3(n7919), .O(n14345) );
  ND2KHD U10400 ( .I1(n10441), .I2(n10091), .O(n7879) );
  ND2KHD U10401 ( .I1(n9832), .I2(n13627), .O(n12404) );
  ND2KHD U10402 ( .I1(n9581), .I2(n12829), .O(n12669) );
  INVGHD U10403 ( .I(n6797), .O(n9260) );
  INVJHD U10404 ( .I(n11802), .O(n7694) );
  INVCKGHD U10405 ( .I(n12781), .O(n8591) );
  ND3EHD U10406 ( .I1(n7112), .I2(n11858), .I3(n7389), .O(n7404) );
  AN2HHD U10407 ( .I1(n11859), .I2(n8886), .O(n7112) );
  ND2HHD U10408 ( .I1(n7113), .I2(n7519), .O(n10267) );
  ND3EHD U10409 ( .I1(n8288), .I2(n9533), .I3(n9535), .O(n7113) );
  ND2HHD U10410 ( .I1(n8167), .I2(n8166), .O(n8165) );
  ND2KHD U10411 ( .I1(n9686), .I2(n10182), .O(n7836) );
  ND2KHD U10412 ( .I1(n9730), .I2(n7864), .O(n8208) );
  BUFEHD U10413 ( .I(n10107), .O(n7114) );
  ND3EHD U10414 ( .I1(n12254), .I2(n11953), .I3(n13409), .O(n11961) );
  NR2GHD U10415 ( .I1(n11950), .I2(n11951), .O(n13409) );
  ND3EHD U10416 ( .I1(n12368), .I2(n13389), .I3(n12369), .O(n12370) );
  ND2HHD U10417 ( .I1(n10098), .I2(n13431), .O(n10097) );
  ND2KHD U10418 ( .I1(n9144), .I2(n12464), .O(n9143) );
  BUFEHD U10419 ( .I(n11508), .O(n7115) );
  ND3EHD U10420 ( .I1(n7333), .I2(n7735), .I3(n12854), .O(n7587) );
  NR2GHD U10421 ( .I1(n10449), .I2(n7734), .O(n7333) );
  ND3EHD U10422 ( .I1(n12728), .I2(n9687), .I3(n12726), .O(n12734) );
  XOR2HHD U10423 ( .I1(n9023), .I2(n9024), .O(n8036) );
  NR2IHD U10424 ( .I1(n8207), .I2(n9444), .O(n10427) );
  NR2EHD U10425 ( .I1(n13437), .I2(n13436), .O(n9058) );
  ND2HHD U10426 ( .I1(n13371), .I2(n9398), .O(n12367) );
  INVGHD U10427 ( .I(n9014), .O(n8111) );
  AN3B1HHD U10428 ( .I1(n9632), .I2(n9216), .B1(n7844), .O(n7843) );
  ND2KHD U10429 ( .I1(n7241), .I2(n7239), .O(n8206) );
  INVNHD U10430 ( .I(n8012), .O(n9694) );
  OAI112BHD U10431 ( .C1(n15503), .C2(n13914), .A1(n7116), .B1(n13921), .O(n6097) );
  ND2HHD U10432 ( .I1(n15503), .I2(n13913), .O(n7116) );
  ND2HHD U10433 ( .I1(n12522), .I2(n8208), .O(n10383) );
  ND2KHD U10434 ( .I1(n8852), .I2(n6901), .O(n7310) );
  ND3EHD U10435 ( .I1(n6641), .I2(n8190), .I3(n11848), .O(n11849) );
  INVNHD U10436 ( .I(n8198), .O(n8199) );
  NR2IHD U10437 ( .I1(n8903), .I2(n11020), .O(n11095) );
  ND3EHD U10438 ( .I1(n8987), .I2(n7878), .I3(n7877), .O(n8885) );
  NR2EHD U10439 ( .I1(n12356), .I2(n12355), .O(n12358) );
  BUFMHD U10440 ( .I(n13053), .O(n7118) );
  ND2HHD U10441 ( .I1(n9397), .I2(n11078), .O(n9704) );
  INVNHD U10442 ( .I(_i_CLEFIA128_keyL _8), .O(n15212) );
  ND2KHD U10443 ( .I1(n7301), .I2(n8188), .O(n12749) );
  ND3EHD U10444 ( .I1(n9873), .I2(n12361), .I3(n12324), .O(n12325) );
  ND3EHD U10445 ( .I1(n14112), .I2(n14110), .I3(n14111), .O(n6203) );
  ND2KHD U10446 ( .I1(n8797), .I2(_i_CLEFIA128_keyK _109), .O(n11889) );
  ND2DHD U10447 ( .I1(n8734), .I2(n7043), .O(n8730) );
  XOR2EHD U10448 ( .I1(n7231), .I2(n14214), .O(n8089) );
  ND3EHD U10449 ( .I1(n7119), .I2(n15073), .I3(_i_CLEFIA128_rndcnt_reg _0), .O(n11887) );
  ND2HHD U10450 ( .I1(n8039), .I2(_i_CLEFIA128_keyK _45), .O(n7119) );
  INVGHD U10451 ( .I(n9619), .O(n8458) );
  INVNHD U10452 ( .I(n7384), .O(n7386) );
  XOR2HHD U10453 ( .I1(n7932), .I2(n9746), .O(n7120) );
  ND3EHD U10454 ( .I1(n6992), .I2(n7122), .I3(n7183), .O(n10861) );
  OR3HHD U10455 ( .I1(n12333), .I2(n9990), .I3(n12434), .O(n7633) );
  ND3EHD U10456 ( .I1(n7496), .I2(n11374), .I3(n12777), .O(n11375) );
  ND2KHD U10457 ( .I1(n12692), .I2(n12867), .O(n9067) );
  ND2HHD U10458 ( .I1(n7126), .I2(n7125), .O(n10542) );
  OR3HHD U10459 ( .I1(n12746), .I2(n7284), .I3(n12565), .O(n7283) );
  ND2KHD U10460 ( .I1(n12226), .I2(n13442), .O(n9342) );
  NR2EHD U10461 ( .I1(n9601), .I2(n10838), .O(n10839) );
  AN2HHD U10462 ( .I1(n13609), .I2(n13608), .O(n13610) );
  MUX2HHD U10463 ( .A(n14217), .B(n14216), .S(n15067), .O(n10010) );
  NR2EHD U10464 ( .I1(n11338), .I2(n11515), .O(n11339) );
  NR2CHD U10465 ( .I1(n7642), .I2(n7127), .O(n11083) );
  NR2IHD U10466 ( .I1(n9187), .I2(n7757), .O(n11997) );
  AN3HHD U10467 ( .I1(n7467), .I2(n7464), .I3(n9603), .O(n8633) );
  ND3EHD U10468 ( .I1(n9463), .I2(n10005), .I3(n7942), .O(n13151) );
  ND3EHD U10469 ( .I1(n8567), .I2(n8566), .I3(n14181), .O(n6162) );
  ND2KHD U10470 ( .I1(n6882), .I2(n9730), .O(n7606) );
  XOR2HHD U10471 ( .I1(DOUT_75), .I2(n8757), .O(n10151) );
  ND3EHD U10472 ( .I1(n7022), .I2(n9310), .I3(n6734), .O(n7749) );
  ND2KHD U10473 ( .I1(n10090), .I2(n8207), .O(n10737) );
  INVGHD U10474 ( .I(n11683), .O(n9043) );
  XOR2KHD U10475 ( .I1(n8400), .I2(n8151), .O(n13216) );
  OAI12CHD U10476 ( .B1(n8519), .B2(n15416), .A1(n14658), .O(n6350) );
  ND3EHD U10477 ( .I1(n10868), .I2(n11078), .I3(n10867), .O(n8900) );
  OA12HHD U10478 ( .B1(n7131), .B2(n9685), .A1(n12591), .O(n9668) );
  ND2KHD U10479 ( .I1(n7133), .I2(n7132), .O(n8181) );
  NR2IHD U10480 ( .I1(n10431), .I2(n8526), .O(n10420) );
  ND2KHD U10481 ( .I1(n9747), .I2(n13590), .O(n12261) );
  ND3EHD U10482 ( .I1(n9125), .I2(n7560), .I3(_i_CLEFIA128_state_reg _1), .O(n7559) );
  ND2KHD U10483 ( .I1(n8899), .I2(_i_CLEFIA128_keyK _44), .O(n9125) );
  NR2EHD U10484 ( .I1(n11643), .I2(n11642), .O(n11645) );
  ND2HHD U10485 ( .I1(n8521), .I2(n8428), .O(n8520) );
  NR2EHD U10486 ( .I1(n12530), .I2(n12540), .O(n11256) );
  OR3HHD U10487 ( .I1(n12627), .I2(n10772), .I3(n10771), .O(n7134) );
  ND3EHD U10488 ( .I1(n7850), .I2(n7849), .I3(n7851), .O(n10017) );
  NR2IHD U10489 ( .I1(n11127), .I2(n11108), .O(n9539) );
  NR2IHD U10490 ( .I1(n10320), .I2(n14707), .O(n10138) );
  BUFMHD U10491 ( .I(n11505), .O(n7546) );
  ND2HHD U10492 ( .I1(n7135), .I2(n9021), .O(n6178) );
  NR2CHD U10493 ( .I1(n8118), .I2(n6981), .O(n7848) );
  ND2HHD U10494 ( .I1(n10092), .I2(n7140), .O(n9819) );
  INVKHD U10495 ( .I(n8176), .O(n7677) );
  ND2KHD U10496 ( .I1(_i_CLEFIA128_keyK _76), .I2(n8797), .O(n7792) );
  ND2KHD U10497 ( .I1(n9209), .I2(n7015), .O(n8801) );
  ND2HHD U10498 ( .I1(n7144), .I2(n7142), .O(n7390) );
  ND2HHD U10499 ( .I1(n11919), .I2(n7143), .O(n7142) );
  OA112EHD U10500 ( .C1(n11915), .C2(n7392), .A1(n7145), .B1(n7391), .O(n7144));
  BUFKHD U10501 ( .I(n11117), .O(n7146) );
  ND3EHD U10502 ( .I1(n7147), .I2(n15277), .I3(_i_CLEFIA128_rndcnt_reg _0), .O(n10319) );
  ND2HHD U10503 ( .I1(n8797), .I2(_i_CLEFIA128_keyK _26), .O(n7147) );
  OA13EHD U10504 ( .B1(n11824), .B2(n11823), .B3(n13075), .A1(n14049), .O(n7148) );
  ND2KHD U10505 ( .I1(n7150), .I2(n7149), .O(n10225) );
  ND3EHD U10506 ( .I1(n7644), .I2(n11587), .I3(n7643), .O(n7149) );
  INVKHD U10507 ( .I(n10419), .O(n10441) );
  ND3EHD U10508 ( .I1(n8557), .I2(n8554), .I3(n8571), .O(n10419) );
  AN3HHD U10509 ( .I1(n7151), .I2(n10872), .I3(n10873), .O(n10880) );
  INVNHD U10510 ( .I(n8205), .O(n8207) );
  OA13EHD U10511 ( .B1(n11481), .B2(n8683), .B3(n11480), .A1(n11479), .O(n11490) );
  ND2HHD U10512 ( .I1(n11028), .I2(n11029), .O(n8683) );
  ND2KHD U10513 ( .I1(n8797), .I2(_i_CLEFIA128_keyK _96), .O(n7557) );
  NR2GHD U10514 ( .I1(n9428), .I2(n9424), .O(n11071) );
  AN3HHD U10515 ( .I1(n13814), .I2(n13844), .I3(n12320), .O(n8718) );
  ND2HHD U10516 ( .I1(n14837), .I2(n15500), .O(n8543) );
  ND2HHD U10517 ( .I1(n10825), .I2(n7052), .O(n8959) );
  NR2CHD U10518 ( .I1(n13831), .I2(n13830), .O(n13832) );
  INVDHD U10519 ( .I(n9672), .O(n11910) );
  ND2KHD U10520 ( .I1(n7163), .I2(n8291), .O(n9672) );
  BUFNHD U10521 ( .I(n10883), .O(n7783) );
  ND3EHD U10522 ( .I1(n8520), .I2(n14324), .I3(n8518), .O(n6099) );
  XNR3EHD U10523 ( .I1(n8486), .I2(n8049), .I3(n14103), .O(n13266) );
  ND3EHD U10524 ( .I1(n11200), .I2(n9598), .I3(n11199), .O(n14103) );
  ND2HHD U10525 ( .I1(n10216), .I2(n6809), .O(n8793) );
  OA12HHD U10526 ( .B1(n7524), .B2(n12840), .A1(n7523), .O(n9622) );
  OR3HHD U10527 ( .I1(n10947), .I2(n10946), .I3(n8909), .O(n8980) );
  ND3CHD U10528 ( .I1(n11114), .I2(n11113), .I3(n11112), .O(n11115) );
  ND3EHD U10529 ( .I1(n11173), .I2(n11457), .I3(n11174), .O(n9599) );
  BUFKHD U10530 ( .I(n8483), .O(n7156) );
  ND2KHD U10531 ( .I1(n12829), .I2(n8215), .O(n10905) );
  NR2GHD U10532 ( .I1(n11623), .I2(n11624), .O(n13492) );
  AN2HHD U10533 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(_i_CLEFIA128_keyL _9), .O(n8380) );
  NR2CHD U10534 ( .I1(n10886), .I2(n7747), .O(n7745) );
  ND2DHD U10535 ( .I1(n7725), .I2(n8295), .O(n10081) );
  ND2HHD U10536 ( .I1(n7329), .I2(n7328), .O(n7327) );
  INVKHD U10537 ( .I(n9579), .O(n9749) );
  NR2GHD U10538 ( .I1(n7344), .I2(n7302), .O(n7157) );
  ND3EHD U10539 ( .I1(n7158), .I2(n8103), .I3(n8104), .O(n7549) );
  ND3EHD U10540 ( .I1(n8109), .I2(n8107), .I3(n8110), .O(n7158) );
  ND3EHD U10541 ( .I1(n8034), .I2(n9420), .I3(n8033), .O(n8032) );
  ND3EHD U10542 ( .I1(n6923), .I2(n12814), .I3(n7753), .O(n7592) );
  NR2GHD U10543 ( .I1(n7749), .I2(n7750), .O(n12814) );
  NR2IHD U10544 ( .I1(_i_CLEFIA128_keyK _64), .I2(n15408), .O(n8108) );
  XNR2KHD U10545 ( .I1(n11975), .I2(n7160), .O(n12001) );
  OAI12CHD U10546 ( .B1(n7814), .B2(n7815), .A1(n12671), .O(n7162) );
  ND2KHD U10547 ( .I1(n9628), .I2(n7335), .O(n13066) );
  NR2IHD U10548 ( .I1(n7720), .I2(n7905), .O(n7825) );
  BUFQHD U10549 ( .I(n10774), .O(n7507) );
  BUFEHD U10550 ( .I(n9774), .O(n7166) );
  ND2HHD U10551 ( .I1(n6805), .I2(n11070), .O(n10359) );
  ND3EHD U10552 ( .I1(n12740), .I2(n8684), .I3(n11029), .O(n7167) );
  NR2GHD U10553 ( .I1(n10663), .I2(n10662), .O(n7168) );
  ND3EHD U10554 ( .I1(n7340), .I2(n8236), .I3(n12867), .O(n8142) );
  OAI112BHD U10555 ( .C1(n14813), .C2(n13987), .A1(n7169), .B1(n13994), .O(n6105) );
  ND2HHD U10556 ( .I1(n14813), .I2(n13986), .O(n7169) );
  ND3EHD U10557 ( .I1(n11974), .I2(n15047), .I3(_i_CLEFIA128_rndcnt_reg _0), .O(n7785) );
  ND2HHD U10558 ( .I1(n7358), .I2(n10267), .O(n7357) );
  ND2HHD U10559 ( .I1(n7875), .I2(n12662), .O(n7358) );
  XOR2HHD U10560 ( .I1(n7170), .I2(n9971), .O(n7577) );
  NR2IHD U10561 ( .I1(n7171), .I2(n12551), .O(n9076) );
  OA12HHD U10562 ( .B1(n9655), .B2(n12527), .A1(n7519), .O(n7171) );
  ND3EHD U10563 ( .I1(n6995), .I2(n9663), .I3(n6671), .O(n12523) );
  ND2HHD U10564 ( .I1(n8521), .I2(n11130), .O(n10041) );
  ND3EHD U10565 ( .I1(n7965), .I2(n12207), .I3(n8795), .O(n9570) );
  XNR3EHD U10566 ( .I1(n14104), .I2(n14245), .I3(n7896), .O(n8091) );
  ND2HHD U10567 ( .I1(n7172), .I2(n10806), .O(n10357) );
  ND2HHD U10568 ( .I1(n7507), .I2(n9730), .O(n7172) );
  OAI112BHD U10569 ( .C1(n6604), .C2(n11129), .A1(n15438), .B1(n7173), .O(n6213) );
  ND2HHD U10570 ( .I1(n15435), .I2(n15500), .O(n7173) );
  XOR2HHD U10571 ( .I1(n7175), .I2(n7174), .O(n15435) );
  XNR3EHD U10572 ( .I1(n14028), .I2(n9768), .I3(n13768), .O(n7174) );
  NR2IHD U10573 ( .I1(n12346), .I2(n7176), .O(n7407) );
  NR2BHD U10574 ( .I1(n7176), .I2(n9875), .O(n9874) );
  INVJHD U10575 ( .I(n9873), .O(n7176) );
  ND3CHD U10576 ( .I1(n10378), .I2(n7178), .I3(n8138), .O(n10379) );
  ND3EHD U10577 ( .I1(n12516), .I2(n7179), .I3(n9656), .O(n9655) );
  ND3EHD U10578 ( .I1(n7179), .I2(n10800), .I3(n10799), .O(n9773) );
  ND3EHD U10579 ( .I1(n11071), .I2(n7179), .I3(n11261), .O(n7875) );
  NR2IHD U10580 ( .I1(n10170), .I2(n10172), .O(n7179) );
  NR2EHD U10581 ( .I1(n10021), .I2(n7181), .O(n9219) );
  INVCKGHD U10582 ( .I(n9211), .O(n7181) );
  AN2KHD U10583 ( .I1(n10324), .I2(n7864), .O(n10021) );
  ND2CHD U10584 ( .I1(n7185), .I2(n7779), .O(n10371) );
  ND2HHD U10585 ( .I1(n12652), .I2(n7185), .O(n11075) );
  ND2HHD U10586 ( .I1(n12623), .I2(n7185), .O(n12653) );
  ND2DHD U10587 ( .I1(n7186), .I2(n11130), .O(n14273) );
  ND2DHD U10588 ( .I1(n7186), .I2(n15500), .O(n14269) );
  ND2DHD U10589 ( .I1(n7186), .I2(n8282), .O(n10078) );
  XNR2KHD U10590 ( .I1(n10063), .I2(n10062), .O(n7186) );
  ND2CHD U10591 ( .I1(n7187), .I2(n9211), .O(n8488) );
  ND2CHD U10592 ( .I1(n7187), .I2(n12623), .O(n10651) );
  ND2KHD U10593 ( .I1(n6842), .I2(n7507), .O(n7187) );
  OR2KHD U10594 ( .I1(n7863), .I2(n9774), .O(n7316) );
  ND2KHD U10595 ( .I1(n7189), .I2(n10660), .O(n9349) );
  AN2HHD U10596 ( .I1(n7188), .I2(n10173), .O(n8889) );
  NR2BHD U10597 ( .I1(n7016), .I2(n9774), .O(n7188) );
  ND2CHD U10598 ( .I1(n7189), .I2(n9766), .O(n10778) );
  OR2EHD U10599 ( .I1(n15513), .I2(n7191), .O(n7211) );
  OAI12CHD U10600 ( .B1(n7191), .B2(n15416), .A1(n14482), .O(n6339) );
  MUX2HHD U10601 ( .A(n13756), .B(n13755), .S(n7191), .O(n13764) );
  XNR3EHD U10602 ( .I1(n13754), .I2(n8766), .I3(n13753), .O(n7191) );
  OR3HHD U10603 ( .I1(n7194), .I2(n7193), .I3(n11064), .O(n11265) );
  XOR2HHD U10604 ( .I1(n8031), .I2(n7195), .O(n14245) );
  AN2HHD U10605 ( .I1(n11484), .I2(n9796), .O(n7196) );
  ND3EHD U10606 ( .I1(n7197), .I2(n10270), .I3(n11088), .O(n9737) );
  ND2HHD U10607 ( .I1(n7198), .I2(n7778), .O(n7774) );
  INVCHD U10608 ( .I(n7776), .O(n7773) );
  OR3HHD U10609 ( .I1(n13576), .I2(n13184), .I3(n7488), .O(n13181) );
  OR3HHD U10610 ( .I1(n8605), .I2(n8706), .I3(n12057), .O(n7488) );
  ND2HHD U10611 ( .I1(n6819), .I2(n11496), .O(n11497) );
  ND2DHD U10612 ( .I1(n6820), .I2(n11510), .O(n7264) );
  ND2KHD U10613 ( .I1(n8116), .I2(n11335), .O(n7200) );
  XOR2HHD U10614 ( .I1(_i_CLEFIA128_keyL _97), .I2(n7202), .O(n11981) );
  ND2HHD U10615 ( .I1(n8797), .I2(_i_CLEFIA128_keyK _97), .O(n7202) );
  OA12HHD U10616 ( .B1(n6899), .B2(n11978), .A1(_i_CLEFIA128_state_reg _1), .O(n7204) );
  ND2HHD U10617 ( .I1(n7205), .I2(n13110), .O(n13108) );
  AN2HHD U10618 ( .I1(n7205), .I2(DOUT_90), .O(n8401) );
  ND2HHD U10619 ( .I1(n8750), .I2(n13622), .O(n7205) );
  ND2KHD U10620 ( .I1(n9050), .I2(n11049), .O(n7206) );
  NR2EHD U10621 ( .I1(n10069), .I2(n6943), .O(n8366) );
  ND2HHD U10622 ( .I1(n9607), .I2(n7028), .O(n11046) );
  OR2CHD U10623 ( .I1(n7029), .I2(n10069), .O(n11040) );
  ND2HHD U10624 ( .I1(n6929), .I2(n7208), .O(n11521) );
  XNR2KHD U10625 ( .I1(n7214), .I2(n7212), .O(n15024) );
  XOR2HHD U10626 ( .I1(n9768), .I2(n14996), .O(n7213) );
  ND2KHD U10627 ( .I1(n11773), .I2(n13643), .O(n13662) );
  ND2KHD U10628 ( .I1(n11681), .I2(n9435), .O(n13643) );
  ND2KHD U10629 ( .I1(n7766), .I2(n10659), .O(n10363) );
  ND2KHD U10630 ( .I1(n7216), .I2(n7215), .O(n7218) );
  NR2GHD U10631 ( .I1(n8199), .I2(n8789), .O(n7215) );
  NR2IHD U10632 ( .I1(n8137), .I2(n10363), .O(n9731) );
  BUFNHD U10633 ( .I(n9731), .O(n7217) );
  INVQHD U10634 ( .I(n7218), .O(n10668) );
  INVCHD U10635 ( .I(n8789), .O(n10173) );
  ND2HHD U10636 ( .I1(n8797), .I2(_i_CLEFIA128_keyK _85), .O(n10556) );
  ND2HHD U10637 ( .I1(n8797), .I2(_i_CLEFIA128_keyK _41), .O(n11881) );
  OR2B1CHD U10638 ( .I1(n8798), .B1(_i_CLEFIA128_keyK _42), .O(n11875) );
  OR2B1CHD U10639 ( .I1(n8798), .B1(_i_CLEFIA128_keyK _19), .O(n10545) );
  ND3EHD U10640 ( .I1(n8797), .I2(n15064), .I3(_i_CLEFIA128_keyK _69), .O(n9791) );
  ND3EHD U10641 ( .I1(n7219), .I2(n14499), .I3(_i_CLEFIA128_keyK _116), .O(n9393) );
  ND3EHD U10642 ( .I1(n8039), .I2(n9502), .I3(_i_CLEFIA128_keyK _125), .O(n11561) );
  ND3EHD U10643 ( .I1(n8797), .I2(n15074), .I3(_i_CLEFIA128_keyK _123), .O(n11576) );
  ND3CHD U10644 ( .I1(n8797), .I2(n15089), .I3(_i_CLEFIA128_keyK _84), .O(n9133) );
  ND3CHD U10645 ( .I1(n7051), .I2(n15069), .I3(_i_CLEFIA128_keyK _81), .O(n10566) );
  ND3EHD U10646 ( .I1(n7221), .I2(n7710), .I3(n6949), .O(n7255) );
  ND3CHD U10647 ( .I1(n7221), .I2(n11054), .I3(n12719), .O(n11055) );
  NR2IHD U10648 ( .I1(n7709), .I2(n7708), .O(n7221) );
  ND2HHD U10649 ( .I1(n7223), .I2(n10964), .O(n10756) );
  ND3CHD U10650 ( .I1(n12832), .I2(n12692), .I3(n7223), .O(n8971) );
  ND2KHD U10651 ( .I1(n8916), .I2(n12829), .O(n7223) );
  ND3EHD U10652 ( .I1(n8947), .I2(n8945), .I3(n8946), .O(n7226) );
  NR2EHD U10653 ( .I1(n10952), .I2(n7229), .O(n7737) );
  ND3EHD U10654 ( .I1(n9735), .I2(n12669), .I3(n12689), .O(n7229) );
  XOR2HHD U10655 ( .I1(n7129), .I2(n7231), .O(n14193) );
  XOR2HHD U10656 ( .I1(n8031), .I2(n8788), .O(n7726) );
  ND2HHD U10657 ( .I1(n7232), .I2(n12671), .O(n8950) );
  ND3EHD U10658 ( .I1(n7768), .I2(n8953), .I3(n8541), .O(n7232) );
  OA13EHD U10659 ( .B1(n10993), .B2(n11545), .B3(n10994), .A1(n12474), .O(n7235) );
  OA13EHD U10660 ( .B1(n10984), .B2(n11467), .B3(n10985), .A1(n12506), .O(n7236) );
  NR2GHD U10661 ( .I1(n7238), .I2(n7237), .O(n8868) );
  OA13EHD U10662 ( .B1(n9919), .B2(n11012), .B3(n11013), .A1(n12462), .O(n7237) );
  OA12HHD U10663 ( .B1(n10184), .B2(n8632), .A1(n12491), .O(n7238) );
  ND2HHD U10664 ( .I1(n7452), .I2(n7240), .O(n7239) );
  AN2HHD U10665 ( .I1(n9448), .I2(n10411), .O(n7240) );
  ND2HHD U10666 ( .I1(n7242), .I2(n9447), .O(n7241) );
  INVQHD U10667 ( .I(_i_CLEFIA128_keyL _12), .O(n14864) );
  ND2CHD U10668 ( .I1(n7243), .I2(n8255), .O(n6336) );
  ND2HHD U10669 ( .I1(n10452), .I2(n7244), .O(n10899) );
  ND2HHD U10670 ( .I1(n8643), .I2(n7245), .O(n13494) );
  ND2HHD U10671 ( .I1(n7245), .I2(n7421), .O(n14068) );
  ND2HHD U10672 ( .I1(n8923), .I2(n10963), .O(n7246) );
  ND2CHD U10673 ( .I1(n7247), .I2(n6647), .O(n10943) );
  ND2KHD U10674 ( .I1(n8916), .I2(n9383), .O(n7247) );
  ND3EHD U10675 ( .I1(_i_CLEFIA128_state_reg _1), .I2(_i_CLEFIA128_keyK _48), .I3(n8797), .O(n7248) );
  ND2HHD U10676 ( .I1(n7250), .I2(_i_CLEFIA128_state_reg _1), .O(n7249) );
  ND2HHD U10677 ( .I1(n7251), .I2(_i_CLEFIA128_rndcnt_reg _0), .O(n7250) );
  XOR2HHD U10678 ( .I1(_i_CLEFIA128_CON_T_x _1), .I2(DOUT_112), .O(n10085));
  OAI112BHD U10679 ( .C1(n15377), .C2(n15513), .A1(n15370), .B1(n15371), .O(n6206) );
  ND3EHD U10680 ( .I1(n7252), .I2(n10900), .I3(n7736), .O(n7445) );
  NR2GHD U10681 ( .I1(n10898), .I2(n7253), .O(n7252) );
  ND3EHD U10682 ( .I1(n12681), .I2(n8564), .I3(n10905), .O(n7253) );
  ND2HHD U10683 ( .I1(n8938), .I2(n7420), .O(n12681) );
  AN2HHD U10684 ( .I1(n9435), .I2(n7254), .O(n12319) );
  NR2IHD U10685 ( .I1(n9830), .I2(n11793), .O(n7930) );
  OA13EHD U10686 ( .B1(n11502), .B2(n7255), .B3(n11501), .A1(n11500), .O(n11519) );
  OA12EHD U10687 ( .B1(n7255), .B2(n8480), .A1(n11479), .O(n7259) );
  ND2KHD U10688 ( .I1(n7042), .I2(n7040), .O(n8095) );
  BUFMHD U10689 ( .I(n9649), .O(n7256) );
  ND3EHD U10690 ( .I1(n7257), .I2(n7260), .I3(n7262), .O(n9649) );
  OA13EHD U10691 ( .B1(n11357), .B2(n8479), .B3(n8683), .A1(n12591), .O(n7258));
  OAI12CHD U10692 ( .B1(n7261), .B2(n9702), .A1(n12575), .O(n7260) );
  OR2EHD U10693 ( .I1(n11055), .I2(n11056), .O(n7261) );
  AO12EHD U10694 ( .B1(n7263), .B2(n8478), .A1(n11044), .O(n7262) );
  ND3EHD U10695 ( .I1(n11933), .I2(n9343), .I3(n7265), .O(n11935) );
  NR2GHD U10696 ( .I1(n12223), .I2(n7266), .O(n7265) );
  ND3EHD U10697 ( .I1(n7269), .I2(n7267), .I3(n12989), .O(n7266) );
  ND3EHD U10698 ( .I1(n8769), .I2(n10986), .I3(n7270), .O(n12507) );
  ND2HHD U10699 ( .I1(n7272), .I2(n12499), .O(n7271) );
  INVCKGHD U10700 ( .I(n12505), .O(n7272) );
  ND2HHD U10701 ( .I1(n11546), .I2(n9136), .O(n12505) );
  ND2HHD U10702 ( .I1(n7276), .I2(n12575), .O(n7275) );
  OR2B1CHD U10703 ( .I1(n12574), .B1(n12569), .O(n7279) );
  ND2HHD U10704 ( .I1(n7281), .I2(n7283), .O(n7280) );
  ND3EHD U10705 ( .I1(n6957), .I2(n7683), .I3(n7496), .O(n7282) );
  OA12HHD U10706 ( .B1(n7287), .B2(n7288), .A1(n12591), .O(n7286) );
  ND3EHD U10707 ( .I1(n7021), .I2(n9025), .I3(n12590), .O(n7287) );
  ND2HHD U10708 ( .I1(n6955), .I2(n12589), .O(n7288) );
  AN2HHD U10709 ( .I1(n7994), .I2(n13826), .O(n7296) );
  OA12HHD U10710 ( .B1(n9484), .B2(n9483), .A1(n14076), .O(n7299) );
  ND2HHD U10711 ( .I1(n8182), .I2(n7301), .O(n11402) );
  ND2HHD U10712 ( .I1(n9898), .I2(n7301), .O(n12585) );
  ND2HHD U10713 ( .I1(n11335), .I2(n7301), .O(n12582) );
  NR2IHD U10714 ( .I1(n6876), .I2(n11504), .O(n7301) );
  OR3HHD U10715 ( .I1(n10331), .I2(n7302), .I3(n10330), .O(n10354) );
  INVCKGHD U10716 ( .I(n7303), .O(n11290) );
  ND2HHD U10717 ( .I1(n12478), .I2(n7304), .O(n7303) );
  ND2HHD U10718 ( .I1(n11552), .I2(n7304), .O(n11005) );
  ND2HHD U10719 ( .I1(n11178), .I2(n7304), .O(n12504) );
  ND2CHD U10720 ( .I1(n12450), .I2(n7304), .O(n11169) );
  ND2KHD U10721 ( .I1(n9087), .I2(n9964), .O(n7304) );
  ND2CHD U10722 ( .I1(n7307), .I2(n12742), .O(n12552) );
  AN2CHD U10723 ( .I1(n7307), .I2(n11382), .O(n7305) );
  AN2CHD U10724 ( .I1(n12558), .I2(n7307), .O(n7306) );
  ND2KHD U10725 ( .I1(n9738), .I2(n9049), .O(n7307) );
  OAI112BHD U10726 ( .C1(n11030), .C2(n11094), .A1(n11503), .B1(n7309), .O(n11031) );
  ND2KHD U10727 ( .I1(n8182), .I2(n8180), .O(n7309) );
  ND2HHD U10728 ( .I1(n12972), .I2(n12973), .O(n13454) );
  ND2KHD U10729 ( .I1(n6639), .I2(n6837), .O(n9806) );
  NR2IHD U10730 ( .I1(n11911), .I2(n9214), .O(n11943) );
  ND3EHD U10731 ( .I1(n14055), .I2(n11644), .I3(n13102), .O(n10156) );
  NR2IHD U10732 ( .I1(n9834), .I2(n9833), .O(n8579) );
  BUFQHD U10733 ( .I(n8226), .O(n8078) );
  ND2KHD U10734 ( .I1(n8078), .I2(n11766), .O(n9605) );
  XNR2KHD U10735 ( .I1(n6577), .I2(n10218), .O(n14332) );
  ND2KHD U10736 ( .I1(n8851), .I2(n9848), .O(n8850) );
  ND2HHD U10737 ( .I1(n14053), .I2(n13066), .O(n8599) );
  ND2KHD U10738 ( .I1(n7292), .I2(n6837), .O(n14072) );
  ND2KHD U10739 ( .I1(n8899), .I2(n8438), .O(n8872) );
  NR2IHD U10740 ( .I1(n7581), .I2(n7582), .O(n9606) );
  NR2CHD U10741 ( .I1(n12921), .I2(n12060), .O(n7960) );
  ND3EHD U10742 ( .I1(n13646), .I2(n12298), .I3(n11813), .O(n11684) );
  ND2HHD U10743 ( .I1(n8797), .I2(_i_CLEFIA128_keyK _74), .O(n10408) );
  ND2KHD U10744 ( .I1(n9581), .I2(n10219), .O(n12796) );
  ND3EHD U10745 ( .I1(n12714), .I2(n12796), .I3(n9003), .O(n10906) );
  ND2KHD U10746 ( .I1(n12030), .I2(n12127), .O(n13208) );
  ND2DHD U10747 ( .I1(n7605), .I2(n8390), .O(n7604) );
  ND3EHD U10748 ( .I1(n8153), .I2(n9207), .I3(n9456), .O(n8871) );
  XNR3EHD U10749 ( .I1(DOUT_20), .I2(n9649), .I3(n10229), .O(n10232) );
  INVJHD U10750 ( .I(n15134), .O(n9595) );
  ND2HHD U10751 ( .I1(n8635), .I2(n9872), .O(n8634) );
  ND2HHD U10752 ( .I1(n8468), .I2(n13268), .O(n8467) );
  NR2GHD U10753 ( .I1(n10024), .I2(n10025), .O(n10022) );
  INVNHD U10754 ( .I(n7310), .O(n10874) );
  OA22EHD U10755 ( .A1(n7166), .A2(n7311), .B1(n9007), .B2(n10637), .O(n12657));
  INVCHD U10756 ( .I(n10874), .O(n7311) );
  ND2KHD U10757 ( .I1(n7312), .I2(n10317), .O(n8986) );
  ND2CHD U10758 ( .I1(n7318), .I2(n10178), .O(n7317) );
  NR2IHD U10759 ( .I1(n10669), .I2(n7024), .O(n7319) );
  ND2HHD U10760 ( .I1(n7323), .I2(n10327), .O(n10355) );
  ND2HHD U10761 ( .I1(n7326), .I2(n7324), .O(n8048) );
  ND2HHD U10762 ( .I1(n7327), .I2(n9949), .O(n7326) );
  NR2IHD U10763 ( .I1(n9951), .I2(n9948), .O(n7329) );
  ND2KHD U10764 ( .I1(n12619), .I2(n6806), .O(n10657) );
  ND2HHD U10765 ( .I1(n7779), .I2(n6805), .O(n10631) );
  ND2HHD U10766 ( .I1(n9344), .I2(n6805), .O(n10843) );
  ND2CHD U10767 ( .I1(n6806), .I2(n12635), .O(n12636) );
  ND2DHD U10768 ( .I1(n11253), .I2(n6805), .O(n10370) );
  ND2KHD U10769 ( .I1(n10802), .I2(n10179), .O(n7330) );
  ND2KHD U10770 ( .I1(n7331), .I2(n10012), .O(n7854) );
  ND2HHD U10771 ( .I1(n8826), .I2(n10309), .O(n7331) );
  NR2IHD U10772 ( .I1(n9943), .I2(n7332), .O(n8826) );
  NR2IHD U10773 ( .I1(n10306), .I2(n14707), .O(n7332) );
  XOR2HHD U10774 ( .I1(n8561), .I2(n13972), .O(n10027) );
  ND2KHD U10775 ( .I1(n7590), .I2(n7585), .O(n8561) );
  ND3EHD U10776 ( .I1(n7821), .I2(n7333), .I3(n9326), .O(n7820) );
  ND2KHD U10777 ( .I1(n9597), .I2(n7335), .O(n13469) );
  ND2KHD U10778 ( .I1(n7034), .I2(n7335), .O(n13096) );
  NR2IHD U10779 ( .I1(n7897), .I2(n11839), .O(n7336) );
  INVCHD U10780 ( .I(n9723), .O(n7341) );
  ND2KHD U10781 ( .I1(n10746), .I2(n9581), .O(n7340) );
  NR2BHD U10782 ( .I1(n9524), .I2(n12836), .O(n10896) );
  NR2EHD U10783 ( .I1(n6925), .I2(n7343), .O(n7978) );
  NR2IHD U10784 ( .I1(n11590), .I2(n14707), .O(n7343) );
  NR2IHD U10785 ( .I1(n7345), .I2(n7346), .O(n12512) );
  ND2KHD U10786 ( .I1(n8797), .I2(_i_CLEFIA128_keyK _77), .O(n7348) );
  ND2HHD U10787 ( .I1(n7349), .I2(n7348), .O(n7351) );
  ND3EHD U10788 ( .I1(n8797), .I2(_i_CLEFIA128_keyK _77), .I3(_i_CLEFIA128_keyL _77), .O(n7350) );
  XOR2HHD U10789 ( .I1(n8088), .I2(n8089), .O(n15095) );
  ND2KHD U10790 ( .I1(n7355), .I2(n7354), .O(n13495) );
  NR2GHD U10791 ( .I1(n9509), .I2(n7027), .O(n7354) );
  ND2HHD U10792 ( .I1(n7359), .I2(n12651), .O(n12628) );
  ND2KHD U10793 ( .I1(n9678), .I2(n7393), .O(n12238) );
  ND2KHD U10794 ( .I1(n11906), .I2(n12226), .O(n9678) );
  ND2KHD U10795 ( .I1(n6905), .I2(n7014), .O(n7361) );
  ND2HHD U10796 ( .I1(n7644), .I2(n7643), .O(n7362) );
  XOR2HHD U10797 ( .I1(n9718), .I2(n7363), .O(n14365) );
  XOR3EHD U10798 ( .I1(DOUT_91), .I2(n7363), .I3(n8755), .O(n8765) );
  ND2KHD U10799 ( .I1(n13160), .I2(n13161), .O(n7363) );
  ND3EHD U10800 ( .I1(n7364), .I2(n12534), .I3(n7018), .O(n12535) );
  ND3EHD U10801 ( .I1(n7364), .I2(n11086), .I3(n8382), .O(n10269) );
  AN2HHD U10802 ( .I1(n9770), .I2(n7954), .O(n13131) );
  ND2KHD U10803 ( .I1(n12125), .I2(n12129), .O(n9770) );
  ND2HHD U10804 ( .I1(n10011), .I2(n9766), .O(n7365) );
  ND3EHD U10805 ( .I1(n9190), .I2(n8193), .I3(n7367), .O(n10947) );
  ND2KHD U10806 ( .I1(n8916), .I2(n10746), .O(n9190) );
  AN2HHD U10807 ( .I1(n9735), .I2(n10945), .O(n7367) );
  AN2HHD U10808 ( .I1(n10905), .I2(n8979), .O(n12704) );
  ND2KHD U10809 ( .I1(n8938), .I2(n10746), .O(n9723) );
  ND2KHD U10810 ( .I1(n8916), .I2(n10219), .O(n12713) );
  NR2GHD U10811 ( .I1(n8740), .I2(n11986), .O(n9318) );
  ND2HHD U10812 ( .I1(n7368), .I2(_i_CLEFIA128_state_reg _1), .O(n8740) );
  ND3EHD U10813 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(n11982), .I3(n15243), .O(n7368) );
  XNR2KHD U10814 ( .I1(_i_CLEFIA128_CON_T_x _2), .I2(DOUT_98), .O(n11986) );
  ND2HHD U10815 ( .I1(n7369), .I2(n13106), .O(n8646) );
  ND2HHD U10816 ( .I1(n12352), .I2(n9093), .O(n13423) );
  ND2KHD U10817 ( .I1(n7037), .I2(n7370), .O(n9093) );
  AN2HHD U10818 ( .I1(n7372), .I2(n7371), .O(n7370) );
  NR2CHD U10819 ( .I1(n8763), .I2(n11911), .O(n7371) );
  NR2CHD U10820 ( .I1(n10209), .I2(n10107), .O(n7372) );
  INVGHD U10821 ( .I(n8453), .O(n12555) );
  ND3EHD U10822 ( .I1(n6954), .I2(n11032), .I3(n7373), .O(n8479) );
  ND2HHD U10823 ( .I1(n10862), .I2(n7375), .O(n9530) );
  ND2HHD U10824 ( .I1(n7375), .I2(n12537), .O(n10782) );
  ND2CHD U10825 ( .I1(n8202), .I2(n7374), .O(n10671) );
  ND2HHD U10826 ( .I1(n7375), .I2(n11253), .O(n12530) );
  ND2CHD U10827 ( .I1(n11067), .I2(n7374), .O(n9428) );
  ND2KHD U10828 ( .I1(n7507), .I2(n10318), .O(n7375) );
  ND3EHD U10829 ( .I1(n9222), .I2(n9031), .I3(n7378), .O(n7377) );
  ND3EHD U10830 ( .I1(n8440), .I2(n10248), .I3(n7379), .O(n10554) );
  ND3EHD U10831 ( .I1(n7380), .I2(n9133), .I3(n7006), .O(n7379) );
  XNR2KHD U10832 ( .I1(n7955), .I2(n9818), .O(n7381) );
  XOR2HHD U10833 ( .I1(n10003), .I2(n7381), .O(n10020) );
  AN2HHD U10834 ( .I1(n7382), .I2(n12268), .O(n12374) );
  ND2HHD U10835 ( .I1(n7382), .I2(n7165), .O(n12035) );
  ND2KHD U10836 ( .I1(n12125), .I2(n8183), .O(n7382) );
  XNR2KHD U10837 ( .I1(n11664), .I2(n7436), .O(n7383) );
  ND2HHD U10838 ( .I1(n11681), .I2(n8200), .O(n10141) );
  INVCKGHD U10839 ( .I(n12349), .O(n11959) );
  ND2KHD U10840 ( .I1(n6823), .I2(n7394), .O(n9516) );
  NR2IHD U10841 ( .I1(n11634), .I2(n11614), .O(n7394) );
  ND2KHD U10842 ( .I1(n7007), .I2(n10005), .O(n7395) );
  NR2IHD U10843 ( .I1(n10848), .I2(n7396), .O(n9146) );
  BUFQHD U10844 ( .I(n11095), .O(n7398) );
  XNR2KHD U10845 ( .I1(n11860), .I2(n7399), .O(n11905) );
  ND2HHD U10846 ( .I1(n7404), .I2(n7400), .O(n7399) );
  NR2GHD U10847 ( .I1(n7402), .I2(n7401), .O(n7400) );
  ND2HHD U10848 ( .I1(n7403), .I2(_i_CLEFIA128_state_reg _1), .O(n7402) );
  ND3EHD U10849 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(n10157), .I3(n15191), .O(n7403) );
  OA13EHD U10850 ( .B1(n7405), .B2(n13363), .B3(n13364), .A1(n13431), .O(n13380) );
  NR2GHD U10851 ( .I1(n12227), .I2(n7406), .O(n10105) );
  NR2GHD U10852 ( .I1(_i_CLEFIA128_keyL _2), .I2(n8589), .O(n8369) );
  INVDHD U10853 ( .I(n9667), .O(n13254) );
  ND2HHD U10854 ( .I1(n7407), .I2(n13000), .O(n11950) );
  AN2HHD U10855 ( .I1(n12432), .I2(n7407), .O(n8402) );
  ND2HHD U10856 ( .I1(n15435), .I2(n11130), .O(n15434) );
  AN2HHD U10857 ( .I1(n7408), .I2(n7858), .O(n12290) );
  NR2GHD U10858 ( .I1(n7409), .I2(n10128), .O(n7858) );
  ND3EHD U10859 ( .I1(n7415), .I2(n7413), .I3(n7411), .O(n7410) );
  ND2HHD U10860 ( .I1(n8576), .I2(n7412), .O(n7411) );
  ND3EHD U10861 ( .I1(n6966), .I2(n8577), .I3(n7414), .O(n7413) );
  ND2HHD U10862 ( .I1(n7416), .I2(n9902), .O(n7415) );
  ND3EHD U10863 ( .I1(n7556), .I2(n6911), .I3(n7867), .O(n12391) );
  ND3CHD U10864 ( .I1(n13581), .I2(n6911), .I3(n13580), .O(n13588) );
  ND2HHD U10865 ( .I1(n7417), .I2(n9998), .O(n12385) );
  AN2CHD U10866 ( .I1(n7417), .I2(n13629), .O(n7552) );
  ND3CHD U10867 ( .I1(n7417), .I2(n13183), .I3(n13595), .O(n12002) );
  ND2KHD U10868 ( .I1(n12125), .I2(n9580), .O(n7417) );
  OA13EHD U10869 ( .B1(n7418), .B2(n11786), .B3(n11785), .A1(n13826), .O(n7583) );
  OA13EHD U10870 ( .B1(n13519), .B2(n13520), .B3(n7418), .A1(n13835), .O(n13536) );
  OR3HHD U10871 ( .I1(n11784), .I2(n11783), .I3(n11782), .O(n7418) );
  OR2KHD U10872 ( .I1(n8760), .I2(n6875), .O(n14043) );
  NR2IHD U10873 ( .I1(n9029), .I2(n9556), .O(n12186) );
  ND2HHD U10874 ( .I1(n13479), .I2(n11644), .O(n12187) );
  ND2KHD U10875 ( .I1(n9597), .I2(n8210), .O(n13479) );
  ND3EHD U10876 ( .I1(n13427), .I2(n12414), .I3(n13430), .O(n7424) );
  ND2HHD U10877 ( .I1(n13448), .I2(n12350), .O(n13375) );
  NR2GHD U10878 ( .I1(n7427), .I2(n13666), .O(n7426) );
  NR2GHD U10879 ( .I1(n12144), .I2(n9815), .O(n8802) );
  ND2HHD U10880 ( .I1(n7432), .I2(n8437), .O(n9982) );
  ND3EHD U10881 ( .I1(n6969), .I2(n10891), .I3(n10890), .O(n7529) );
  ND3EHD U10882 ( .I1(n6969), .I2(n9963), .I3(n10757), .O(n10827) );
  NR2GHD U10883 ( .I1(n9419), .I2(n8498), .O(n8034) );
  ND2HHD U10884 ( .I1(n7435), .I2(_i_CLEFIA128_state_reg _1), .O(n9419) );
  XNR2HHD U10885 ( .I1(_i_CLEFIA128_CON_T_x _9), .I2(DOUT_56), .O(n8498) );
  ND2HHD U10886 ( .I1(n7438), .I2(n7437), .O(n9495) );
  ND3EHD U10887 ( .I1(n13851), .I2(n13850), .I3(DOUT_92), .O(n7437) );
  ND2HHD U10888 ( .I1(n7439), .I2(n9496), .O(n7438) );
  NR2IHD U10889 ( .I1(n8053), .I2(n8055), .O(n13850) );
  ND2CHD U10890 ( .I1(n7931), .I2(n7440), .O(n12082) );
  ND2HHD U10891 ( .I1(n12296), .I2(n7440), .O(n7786) );
  ND3EHD U10892 ( .I1(n7931), .I2(n9621), .I3(n7440), .O(n13654) );
  ND2KHD U10893 ( .I1(n6872), .I2(n7386), .O(n7440) );
  ND2HHD U10894 ( .I1(n13401), .I2(n12366), .O(n7441) );
  XOR2HHD U10895 ( .I1(n7836), .I2(n10217), .O(n14331) );
  XNR3EHD U10896 ( .I1(n14345), .I2(n13556), .I3(n7836), .O(n8988) );
  XNR3EHD U10897 ( .I1(DOUT_83), .I2(n8578), .I3(n7836), .O(n14363) );
  NR2CHD U10898 ( .I1(n12413), .I2(n7442), .O(n11944) );
  ND3EHD U10899 ( .I1(n8289), .I2(n13421), .I3(n13460), .O(n7442) );
  ND2HHD U10900 ( .I1(n7443), .I2(n8529), .O(n7523) );
  ND3EHD U10901 ( .I1(n12783), .I2(n8352), .I3(n10903), .O(n7446) );
  ND2HHD U10902 ( .I1(n6976), .I2(n7737), .O(n7447) );
  ND2HHD U10903 ( .I1(n7450), .I2(n8758), .O(n7941) );
  ND2CHD U10904 ( .I1(n7450), .I2(n12320), .O(n11815) );
  AN2HHD U10905 ( .I1(n7450), .I2(n13642), .O(n8610) );
  ND2HHD U10906 ( .I1(n11709), .I2(n7450), .O(n11710) );
  AN2CHD U10907 ( .I1(n12092), .I2(n6682), .O(n7449) );
  ND2KHD U10908 ( .I1(n9811), .I2(n7035), .O(n7450) );
  NR2GHD U10909 ( .I1(n8437), .I2(n9771), .O(n8825) );
  ND3EHD U10910 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(n11962), .I3(n15182), .O(n7453) );
  XNR2HHD U10911 ( .I1(_i_CLEFIA128_CON_T_xi_2 ), .I2(DOUT_100), .O(n8437) );
  INVJHD U10912 ( .I(n7454), .O(n10450) );
  ND2KHD U10913 ( .I1(n8908), .I2(n12829), .O(n7454) );
  ND2HHD U10914 ( .I1(n7454), .I2(n10755), .O(n8917) );
  ND2HHD U10915 ( .I1(n8914), .I2(n7456), .O(n8913) );
  AN2HHD U10916 ( .I1(n9095), .I2(n6938), .O(n9044) );
  ND3EHD U10917 ( .I1(n7533), .I2(n7534), .I3(n11676), .O(n7458) );
  ND3EHD U10918 ( .I1(n7464), .I2(n7460), .I3(n9603), .O(n7459) );
  ND2HHD U10919 ( .I1(n7470), .I2(n7467), .O(n7461) );
  ND3EHD U10920 ( .I1(n7462), .I2(n10134), .I3(n12290), .O(n9882) );
  NR2EHD U10921 ( .I1(n7463), .I2(n13576), .O(n7470) );
  ND2HHD U10922 ( .I1(n15207), .I2(n11130), .O(n8602) );
  XNR2KHD U10923 ( .I1(n13961), .I2(n7471), .O(n15207) );
  XOR2HHD U10924 ( .I1(n14490), .I2(n7724), .O(n8910) );
  ND2KHD U10925 ( .I1(n9622), .I2(n10216), .O(n7724) );
  XOR2HHD U10926 ( .I1(DOUT_15), .I2(n14489), .O(n7472) );
  ND2KHD U10927 ( .I1(n9782), .I2(n9783), .O(n14489) );
  ND2HHD U10928 ( .I1(n8338), .I2(n7473), .O(n11328) );
  ND2HHD U10929 ( .I1(n6817), .I2(n8470), .O(n8004) );
  INVNHD U10930 ( .I(n9327), .O(n9559) );
  ND2HHD U10931 ( .I1(n12681), .I2(n10899), .O(n12789) );
  ND2HHD U10932 ( .I1(n7475), .I2(n8511), .O(n12791) );
  OR3HHD U10933 ( .I1(n7649), .I2(n8882), .I3(n7478), .O(n7480) );
  NR2IHD U10934 ( .I1(n7482), .I2(n7483), .O(n7481) );
  NR2IHD U10935 ( .I1(n10458), .I2(n14707), .O(n7483) );
  OA13CHD U10936 ( .B1(n13378), .B2(n13377), .B3(n7484), .A1(n8264), .O(n13379) );
  OA13EHD U10937 ( .B1(n7485), .B2(n10368), .B3(n10367), .A1(n7519), .O(n7600));
  OA13EHD U10938 ( .B1(n7485), .B2(n12664), .B3(n12663), .A1(n12662), .O(n9308) );
  OA13EHD U10939 ( .B1(n12632), .B2(n12649), .B3(n7485), .A1(n7519), .O(n9305));
  ND3EHD U10940 ( .I1(n10361), .I2(n10360), .I3(n9457), .O(n7485) );
  ND2KHD U10941 ( .I1(n9084), .I2(n7487), .O(n12967) );
  ND2HHD U10942 ( .I1(n7487), .I2(n13439), .O(n12240) );
  ND2CHD U10943 ( .I1(n7487), .I2(n9225), .O(n9608) );
  ND2HHD U10944 ( .I1(n13458), .I2(n7486), .O(n13463) );
  ND3HHD U10945 ( .I1(n13441), .I2(n9679), .I3(n7486), .O(n11958) );
  ND2KHD U10946 ( .I1(n12424), .I2(n7032), .O(n7487) );
  INVCKGHD U10947 ( .I(n12749), .O(n7492) );
  OA13EHD U10948 ( .B1(n11361), .B2(n7494), .B3(n11362), .A1(n11500), .O(n9724) );
  ND3EHD U10949 ( .I1(n8474), .I2(n11342), .I3(n6948), .O(n11362) );
  ND3CHD U10950 ( .I1(n7496), .I2(n11123), .I3(n7115), .O(n11124) );
  NR2IHD U10951 ( .I1(n11118), .I2(n7685), .O(n7496) );
  ND2HHD U10952 ( .I1(n7499), .I2(n11506), .O(n11111) );
  ND2KHD U10953 ( .I1(n8116), .I2(n9801), .O(n7499) );
  OR3HHD U10954 ( .I1(n13244), .I2(n7502), .I3(n9892), .O(n14069) );
  ND2HHD U10955 ( .I1(n13085), .I2(n13469), .O(n7502) );
  ND2KHD U10956 ( .I1(n10095), .I2(n9580), .O(n13572) );
  ND2KHD U10957 ( .I1(n12900), .I2(n12127), .O(n12123) );
  NR2IHD U10958 ( .I1(n9330), .I2(n12520), .O(n10774) );
  ND2HHD U10959 ( .I1(n7510), .I2(n13634), .O(n7509) );
  ND3EHD U10960 ( .I1(n8363), .I2(n7511), .I3(n8633), .O(n7510) );
  ND2HHD U10961 ( .I1(n7513), .I2(n13585), .O(n7512) );
  OR3HHD U10962 ( .I1(n13635), .I2(n12286), .I3(n13169), .O(n7513) );
  AN2HHD U10963 ( .I1(n7516), .I2(n7515), .O(n7514) );
  OAI12CHD U10964 ( .B1(n12275), .B2(n7957), .A1(n13608), .O(n7515) );
  ND3EHD U10965 ( .I1(n7961), .I2(n12061), .I3(n7960), .O(n12275) );
  OAI13BHD U10966 ( .B1(n7518), .B2(n7517), .B3(n10033), .A1(n13622), .O(n7516) );
  ND3EHD U10967 ( .I1(n12389), .I2(n12263), .I3(n12274), .O(n10033) );
  ND3EHD U10968 ( .I1(n12259), .I2(n12923), .I3(n12257), .O(n7517) );
  ND3EHD U10969 ( .I1(n12258), .I2(n12270), .I3(n12269), .O(n7518) );
  ND2HHD U10970 ( .I1(n6803), .I2(n11230), .O(n11087) );
  ND2HHD U10971 ( .I1(n7520), .I2(n8975), .O(n8942) );
  ND2KHD U10972 ( .I1(n8899), .I2(n8317), .O(n8943) );
  INVQHD U10973 ( .I(n14707), .O(n8899) );
  ND2HHD U10974 ( .I1(n9378), .I2(n10895), .O(n7526) );
  NR2IHD U10975 ( .I1(n7528), .I2(n7527), .O(n10216) );
  OA12HHD U10976 ( .B1(n8937), .B2(n10887), .A1(n10282), .O(n7527) );
  ND2HHD U10977 ( .I1(n9939), .I2(n8359), .O(n8937) );
  OA13EHD U10978 ( .B1(n7529), .B2(n10892), .B3(n12667), .A1(n12671), .O(n7528) );
  ND2HHD U10979 ( .I1(n7794), .I2(n8494), .O(n10892) );
  ND2HHD U10980 ( .I1(n10341), .I2(n7530), .O(n10342) );
  OA12HHD U10981 ( .B1(n10336), .B2(_i_CLEFIA128_keyL _94), .A1(n7531), .O(n7530) );
  OAI12CHD U10982 ( .B1(n7578), .B2(n11674), .A1(n8310), .O(n7533) );
  ND3EHD U10983 ( .I1(n7535), .I2(n10148), .I3(n7536), .O(n7534) );
  NR2GHD U10984 ( .I1(n8310), .I2(n11674), .O(n7535) );
  ND2HHD U10985 ( .I1(n7537), .I2(n13642), .O(n7787) );
  ND2CHD U10986 ( .I1(n7537), .I2(n13838), .O(n13840) );
  ND2KHD U10987 ( .I1(n9807), .I2(n8209), .O(n7537) );
  BUFGHD U10988 ( .I(n12172), .O(n7538) );
  ND2KHD U10989 ( .I1(n12172), .I2(n7808), .O(n8292) );
  AN2HHD U10990 ( .I1(n12737), .I2(n7539), .O(n10535) );
  ND2KHD U10991 ( .I1(n8182), .I2(n11049), .O(n7539) );
  ND2HHD U10992 ( .I1(n8663), .I2(n7541), .O(n7540) );
  ND2KHD U10993 ( .I1(n8797), .I2(_i_CLEFIA128_keyK _117), .O(n11661) );
  INVGHD U10994 ( .I(_i_CLEFIA128_keyL _117), .O(n7544) );
  ND2HHD U10995 ( .I1(n7542), .I2(_i_CLEFIA128_state_reg _1), .O(n7989) );
  ND2HHD U10996 ( .I1(n7545), .I2(n7543), .O(n7542) );
  NR2GHD U10997 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(n7544), .O(n7543) );
  INVKHD U10998 ( .I(n7550), .O(n8175) );
  ND2HHD U10999 ( .I1(n8175), .I2(n7031), .O(n7551) );
  ND2KHD U11000 ( .I1(n12125), .I2(n12127), .O(n13596) );
  ND2HHD U11001 ( .I1(n13602), .I2(n12287), .O(n12388) );
  ND2KHD U11002 ( .I1(n12900), .I2(n8183), .O(n8657) );
  ND2KHD U11003 ( .I1(n12291), .I2(n13132), .O(n12402) );
  ND2HHD U11004 ( .I1(n8135), .I2(n7010), .O(n13126) );
  XOR2HHD U11005 ( .I1(_i_CLEFIA128_keyL _96), .I2(n7557), .O(n11990) );
  ND2KHD U11006 ( .I1(n7558), .I2(n9267), .O(n9266) );
  ND2HHD U11007 ( .I1(n7565), .I2(n7563), .O(n7562) );
  NR2GHD U11008 ( .I1(n7564), .I2(n12238), .O(n7563) );
  ND2HHD U11009 ( .I1(n13444), .I2(n9093), .O(n7564) );
  ND3EHD U11010 ( .I1(n13005), .I2(n13028), .I3(n13399), .O(n12237) );
  ND2KHD U11011 ( .I1(n8797), .I2(_i_CLEFIA128_keyK _3), .O(n7566) );
  OR3HHD U11012 ( .I1(n11494), .I2(n9036), .I3(n10515), .O(n11038) );
  ND2HHD U11013 ( .I1(n7568), .I2(_i_CLEFIA128_keyK _67), .O(n8019) );
  NR2GHD U11014 ( .I1(n8798), .I2(_i_CLEFIA128_keyL _67), .O(n7568) );
  OAI112BHD U11015 ( .C1(n10076), .C2(n14353), .A1(n7569), .B1(n14360), .O(n6148) );
  ND2KHD U11016 ( .I1(n10076), .I2(n8261), .O(n7569) );
  XNR2KHD U11017 ( .I1(n7573), .I2(n7570), .O(n10076) );
  XOR2HHD U11018 ( .I1(n7572), .I2(n7571), .O(n7570) );
  XOR2HHD U11019 ( .I1(n10149), .I2(n14352), .O(n7571) );
  XOR2HHD U11020 ( .I1(n14635), .I2(n8830), .O(n7573) );
  ND2CHD U11021 ( .I1(n11699), .I2(n6843), .O(n11701) );
  ND2CHD U11022 ( .I1(n11689), .I2(n6843), .O(n11691) );
  ND2CHD U11023 ( .I1(n10402), .I2(n6843), .O(n10404) );
  ND2CHD U11024 ( .I1(n11917), .I2(n6843), .O(n11919) );
  ND2CHD U11025 ( .I1(n10576), .I2(n6843), .O(n10578) );
  ND2CHD U11026 ( .I1(n12018), .I2(n6843), .O(n12020) );
  ND2HHD U11027 ( .I1(n7574), .I2(n11605), .O(n11607) );
  ND2CHD U11028 ( .I1(n10392), .I2(n6843), .O(n10394) );
  ND2CHD U11029 ( .I1(n12010), .I2(n6843), .O(n12012) );
  ND2CHD U11030 ( .I1(n10500), .I2(n6843), .O(n10501) );
  ND2CHD U11031 ( .I1(n10490), .I2(n6843), .O(n10492) );
  ND2CHD U11032 ( .I1(n10604), .I2(n6843), .O(n10606) );
  ND2KHD U11033 ( .I1(n10337), .I2(n8798), .O(n7574) );
  ND2KHD U11034 ( .I1(n12190), .I2(n7292), .O(n9185) );
  XOR2HHD U11035 ( .I1(n7577), .I2(n9550), .O(n10231) );
  XOR2HHD U11036 ( .I1(n7577), .I2(n9756), .O(n13973) );
  XNR3EHD U11037 ( .I1(n12886), .I2(n7577), .I3(n8651), .O(n10062) );
  OA12HHD U11038 ( .B1(n8819), .B2(n8817), .A1(n8294), .O(n7581) );
  OA12HHD U11039 ( .B1(n8835), .B2(n8837), .A1(n13835), .O(n7584) );
  ND2HHD U11040 ( .I1(n7587), .I2(n9872), .O(n7586) );
  ND2HHD U11041 ( .I1(n7589), .I2(n12671), .O(n7588) );
  OA112HHD U11042 ( .C1(n7719), .C2(n8562), .A1(n7591), .B1(n8528), .O(n7590));
  ND2HHD U11043 ( .I1(n7592), .I2(n10282), .O(n7591) );
  ND2HHD U11044 ( .I1(n14046), .I2(n7594), .O(n7593) );
  ND2HHD U11045 ( .I1(n7595), .I2(n13526), .O(n8836) );
  ND3EHD U11046 ( .I1(n7595), .I2(n8840), .I3(n13819), .O(n12074) );
  NR2GHD U11047 ( .I1(n8834), .I2(n9217), .O(n7595) );
  ND2HHD U11048 ( .I1(n7783), .I2(n8133), .O(n7596) );
  OA13EHD U11049 ( .B1(n10355), .B2(n10354), .B3(n12648), .A1(n12646), .O(n7599) );
  OR2HHD U11050 ( .I1(n7603), .I2(n7605), .O(n8544) );
  OR2HHD U11051 ( .I1(n15513), .I2(n7605), .O(n8567) );
  XOR2HHD U11052 ( .I1(n10196), .I2(n10195), .O(n7605) );
  ND2HHD U11053 ( .I1(n7606), .I2(n8235), .O(n10658) );
  AN2HHD U11054 ( .I1(n12652), .I2(n7606), .O(n8040) );
  XNR3EHD U11055 ( .I1(n8486), .I2(n7607), .I3(n9415), .O(n14244) );
  ND2KHD U11056 ( .I1(n10268), .I2(n8030), .O(n7607) );
  OAI12CHD U11057 ( .B1(n9156), .B2(n7611), .A1(n10181), .O(n9986) );
  ND2HHD U11058 ( .I1(n7609), .I2(n13835), .O(n7923) );
  ND3EHD U11059 ( .I1(n7925), .I2(n6963), .I3(n7926), .O(n7609) );
  ND2HHD U11060 ( .I1(n7610), .I2(n8294), .O(n7922) );
  OR3HHD U11061 ( .I1(n7873), .I2(n13848), .I3(n13849), .O(n7610) );
  INVCKGHD U11062 ( .I(n14343), .O(n7611) );
  ND2KHD U11063 ( .I1(n7612), .I2(n13817), .O(n14343) );
  ND3EHD U11064 ( .I1(n7846), .I2(n7845), .I3(n6965), .O(n7612) );
  ND2KHD U11065 ( .I1(n9042), .I2(n8199), .O(n9562) );
  MUX2HHD U11066 ( .A(n14248), .B(n14247), .S(n8074), .O(n8163) );
  OR3HHD U11067 ( .I1(n11684), .I2(n7938), .I3(n8848), .O(n13666) );
  ND2HHD U11068 ( .I1(n8333), .I2(n12303), .O(n7614) );
  ND2KHD U11069 ( .I1(n7617), .I2(n10290), .O(n13264) );
  ND2DHD U11070 ( .I1(n7617), .I2(n7043), .O(n7616) );
  XNR2KHD U11071 ( .I1(n10117), .I2(n10116), .O(n7617) );
  AN2HHD U11072 ( .I1(n9593), .I2(n7900), .O(n12473) );
  ND2KHD U11073 ( .I1(n10600), .I2(n8767), .O(n7900) );
  ND3EHD U11074 ( .I1(n10235), .I2(n13429), .I3(n9301), .O(n7632) );
  ND3EHD U11075 ( .I1(n7622), .I2(n7631), .I3(n7630), .O(n13215) );
  ND2HHD U11076 ( .I1(n7625), .I2(n7624), .O(n7623) );
  ND2HHD U11077 ( .I1(n11935), .I2(n8264), .O(n7624) );
  ND2HHD U11078 ( .I1(n11927), .I2(n13458), .O(n7625) );
  ND3EHD U11079 ( .I1(n7628), .I2(n7629), .I3(n7627), .O(n7626) );
  ND2HHD U11080 ( .I1(n13381), .I2(n6939), .O(n7627) );
  ND2HHD U11081 ( .I1(n11926), .I2(n13458), .O(n7629) );
  XOR2HHD U11082 ( .I1(n12373), .I2(n13215), .O(n9519) );
  OAI12CHD U11083 ( .B1(n11946), .B2(n11945), .A1(n13431), .O(n7630) );
  ND2HHD U11084 ( .I1(n7635), .I2(n8264), .O(n7634) );
  ND3EHD U11085 ( .I1(n12358), .I2(n9221), .I3(n12357), .O(n7635) );
  ND2HHD U11086 ( .I1(n7637), .I2(n13426), .O(n7636) );
  ND3EHD U11087 ( .I1(n12372), .I2(n9301), .I3(n9117), .O(n7637) );
  ND2KHD U11088 ( .I1(n10720), .I2(n7639), .O(n10972) );
  ND2KHD U11089 ( .I1(n7641), .I2(n10051), .O(n8177) );
  INVCKIHD U11090 ( .I(n7698), .O(n7697) );
  ND2HHD U11091 ( .I1(n9300), .I2(n13651), .O(n7698) );
  NR2IHD U11092 ( .I1(n9890), .I2(n9891), .O(n7644) );
  ND2KHD U11093 ( .I1(n9186), .I2(n11766), .O(n13078) );
  ND3EHD U11094 ( .I1(n6933), .I2(n13078), .I3(n13217), .O(n9357) );
  BUFGHD U11095 ( .I(n10228), .O(n7648) );
  NR2GHD U11096 ( .I1(n7648), .I2(n8897), .O(n12031) );
  ND2HHD U11097 ( .I1(n9777), .I2(n7648), .O(n10130) );
  ND2HHD U11098 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(_i_CLEFIA128_keyL _3), .O(n7654) );
  INVGHD U11099 ( .I(n8015), .O(n11413) );
  NR2GHD U11100 ( .I1(n11089), .I2(n11395), .O(n11322) );
  NR2GHD U11101 ( .I1(n6896), .I2(n11111), .O(n7656) );
  AN2HHD U11102 ( .I1(n7657), .I2(n12577), .O(n11098) );
  ND2HHD U11103 ( .I1(n6789), .I2(n9607), .O(n10538) );
  ND2KHD U11104 ( .I1(n8116), .I2(n8182), .O(n7657) );
  ND2HHD U11105 ( .I1(n7658), .I2(n12575), .O(n7663) );
  ND3EHD U11106 ( .I1(n7662), .I2(n11413), .I3(n6953), .O(n7661) );
  ND2HHD U11107 ( .I1(n11407), .I2(n11404), .O(n7665) );
  ND2HHD U11108 ( .I1(n12091), .I2(n7669), .O(n8620) );
  ND2KHD U11109 ( .I1(n7671), .I2(n7621), .O(n9531) );
  ND2HHD U11110 ( .I1(n10281), .I2(n10587), .O(n11547) );
  ND3EHD U11111 ( .I1(n10513), .I2(n12586), .I3(n7673), .O(n10514) );
  ND3EHD U11112 ( .I1(n8373), .I2(n9687), .I3(n7673), .O(n11381) );
  INVCKGHD U11113 ( .I(n7675), .O(n12770) );
  NR2GHD U11114 ( .I1(n7014), .I2(n8176), .O(n7675) );
  ND2HHD U11115 ( .I1(n7679), .I2(n12563), .O(n7678) );
  ND3EHD U11116 ( .I1(n9682), .I2(n12752), .I3(n12564), .O(n7684) );
  ND2HHD U11117 ( .I1(n7688), .I2(n7691), .O(n10056) );
  ND2HHD U11118 ( .I1(n6959), .I2(n7696), .O(n7690) );
  AN3HHD U11119 ( .I1(n7693), .I2(n12301), .I3(n7692), .O(n7691) );
  ND2HHD U11120 ( .I1(n6912), .I2(n7696), .O(n13675) );
  ND2HHD U11121 ( .I1(n7697), .I2(n12320), .O(n11803) );
  ND3EHD U11122 ( .I1(n10187), .I2(n7699), .I3(n11574), .O(n8022) );
  NR2IHD U11123 ( .I1(n10189), .I2(n10190), .O(n7699) );
  ND2KHD U11124 ( .I1(n8655), .I2(n13810), .O(n7700) );
  INVCKGHD U11125 ( .I(n12143), .O(n7701) );
  NR2EHD U11126 ( .I1(n7700), .I2(n13532), .O(n8614) );
  NR2GHD U11127 ( .I1(n9813), .I2(n7700), .O(n9812) );
  NR2BHD U11128 ( .I1(n7700), .I2(n12305), .O(n10035) );
  ND2HHD U11129 ( .I1(n6837), .I2(n7704), .O(n9511) );
  INVCHD U11130 ( .I(n12189), .O(n7704) );
  BUFGHD U11131 ( .I(n11402), .O(n7705) );
  NR2GHD U11132 ( .I1(n7707), .I2(n9340), .O(n13823) );
  ND2HHD U11133 ( .I1(n9612), .I2(n13804), .O(n9340) );
  INVCKGHD U11134 ( .I(n13837), .O(n7707) );
  ND3EHD U11135 ( .I1(n12727), .I2(n11340), .I3(n11403), .O(n7708) );
  ND2KHD U11136 ( .I1(n11335), .I2(n12561), .O(n11403) );
  INVLHD U11137 ( .I(_i_CLEFIA128_keyL _69), .O(n15064) );
  OA13EHD U11138 ( .B1(n8828), .B2(n14088), .B3(n14089), .A1(n14087), .O(n7711) );
  ND2HHD U11139 ( .I1(n6742), .I2(n7714), .O(n7713) );
  ND2HHD U11140 ( .I1(n15481), .I2(n11130), .O(n14771) );
  XOR2HHD U11141 ( .I1(n14768), .I2(n7715), .O(n15481) );
  XOR2HHD U11142 ( .I1(n9362), .I2(n14767), .O(n7715) );
  XOR2HHD U11143 ( .I1(n8746), .I2(n9816), .O(n14767) );
  XNR2KHD U11144 ( .I1(n10409), .I2(n7727), .O(n7721) );
  ND2HHD U11145 ( .I1(n10883), .I2(n7721), .O(n10938) );
  ND2HHD U11146 ( .I1(n7721), .I2(n10446), .O(n10426) );
  NR2GHD U11147 ( .I1(n7720), .I2(n10755), .O(n9059) );
  NR2IHD U11148 ( .I1(n12703), .I2(n8964), .O(n7751) );
  ND2KHD U11149 ( .I1(n7722), .I2(n8888), .O(n12703) );
  XOR2HHD U11150 ( .I1(n7724), .I2(n9971), .O(n8719) );
  ND2DHD U11151 ( .I1(n7725), .I2(n15500), .O(n14179) );
  ND2DHD U11152 ( .I1(n7725), .I2(n7043), .O(n10174) );
  OA12HHD U11153 ( .B1(n7725), .B2(n14258), .A1(n14265), .O(n10082) );
  XNR2KHD U11154 ( .I1(n10211), .I2(n10083), .O(n7725) );
  XOR2HHD U11155 ( .I1(n10027), .I2(n7726), .O(n8981) );
  ND3EHD U11156 ( .I1(n7033), .I2(n8565), .I3(n8615), .O(n7731) );
  ND2HHD U11157 ( .I1(n12797), .I2(n10759), .O(n7728) );
  ND3EHD U11158 ( .I1(n6915), .I2(n6916), .I3(n9190), .O(n7734) );
  NR2IHD U11159 ( .I1(n8931), .I2(n8934), .O(n10891) );
  INVCKGHD U11160 ( .I(n8917), .O(n7736) );
  ND2HHD U11161 ( .I1(n10960), .I2(n8914), .O(n10952) );
  ND3EHD U11162 ( .I1(n7741), .I2(n12885), .I3(n7738), .O(n14169) );
  ND2HHD U11163 ( .I1(n7739), .I2(n10282), .O(n7738) );
  ND2HHD U11164 ( .I1(n6974), .I2(n7740), .O(n7739) );
  AN2HHD U11165 ( .I1(n12853), .I2(n12854), .O(n7743) );
  OR2EHD U11166 ( .I1(n12874), .I2(n12875), .O(n12882) );
  ND2KHD U11167 ( .I1(n8236), .I2(n12790), .O(n12874) );
  ND2KHD U11168 ( .I1(n7825), .I2(n10123), .O(n8236) );
  ND2KHD U11169 ( .I1(n8859), .I2(n7744), .O(n9644) );
  INVJHD U11170 ( .I(n7783), .O(n7744) );
  ND2HHD U11171 ( .I1(n6968), .I2(n7746), .O(n12680) );
  NR2GHD U11172 ( .I1(n10735), .I2(n12683), .O(n7753) );
  ND2HHD U11173 ( .I1(n6971), .I2(n10810), .O(n12683) );
  ND2KHD U11174 ( .I1(n8240), .I2(n8377), .O(n10735) );
  ND2KHD U11175 ( .I1(n9723), .I2(n12847), .O(n8965) );
  INVGHD U11176 ( .I(n7755), .O(n7752) );
  ND2HHD U11177 ( .I1(n8962), .I2(n12688), .O(n7755) );
  INVCKGHD U11178 ( .I(n9310), .O(n7754) );
  OR3HHD U11179 ( .I1(n7755), .I2(n8970), .I3(n7754), .O(n9302) );
  ND2HHD U11180 ( .I1(n7752), .I2(n7751), .O(n7750) );
  ND2HHD U11181 ( .I1(n8411), .I2(n7783), .O(n7756) );
  NR2IHD U11182 ( .I1(n6881), .I2(n7757), .O(n12004) );
  ND2KHD U11183 ( .I1(n12914), .I2(n10228), .O(n7757) );
  ND2KHD U11184 ( .I1(n7758), .I2(n8077), .O(n9565) );
  OA12HHD U11185 ( .B1(n7760), .B2(n7761), .A1(n7763), .O(n9566) );
  NR2IHD U11186 ( .I1(n11567), .I2(n6741), .O(n7760) );
  ND2DHD U11187 ( .I1(n11569), .I2(_i_CLEFIA128_state_reg _1), .O(n7761) );
  OR3HHD U11188 ( .I1(n13253), .I2(n13254), .I3(n13472), .O(n7764) );
  ND2HHD U11189 ( .I1(n7765), .I2(n9947), .O(n9865) );
  OA13EHD U11190 ( .B1(n13454), .B2(n12974), .B3(n8625), .A1(n13426), .O(n9946) );
  OA12HHD U11191 ( .B1(n12960), .B2(n12961), .A1(n13431), .O(n9945) );
  INVCHD U11192 ( .I(n7034), .O(n13219) );
  ND2HHD U11193 ( .I1(n13182), .I2(n12376), .O(n12400) );
  ND2KHD U11194 ( .I1(n7766), .I2(n10325), .O(n10332) );
  ND3EHD U11195 ( .I1(n10954), .I2(n10955), .I3(n10953), .O(n7767) );
  ND2HHD U11196 ( .I1(n8957), .I2(n9872), .O(n7770) );
  ND2HHD U11197 ( .I1(n8980), .I2(n10282), .O(n7771) );
  ND2HHD U11198 ( .I1(n8955), .I2(n10282), .O(n7772) );
  XNR2KHD U11199 ( .I1(_i_CLEFIA128_CON_T_xi_2 ), .I2(DOUT_115), .O(n9175) );
  ND2HHD U11200 ( .I1(n8168), .I2(n8169), .O(n6209) );
  ND2HHD U11201 ( .I1(n7779), .I2(n11070), .O(n10863) );
  ND2CHD U11202 ( .I1(n7779), .I2(n12609), .O(n12525) );
  ND2KHD U11203 ( .I1(n9730), .I2(n10668), .O(n7779) );
  AN2HHD U11204 ( .I1(n8587), .I2(_i_CLEFIA128_state_reg _1), .O(n7782) );
  ND3EHD U11205 ( .I1(n8942), .I2(n8939), .I3(n8972), .O(n10883) );
  OA112HHD U11206 ( .C1(n11974), .C2(n11973), .A1(n7785), .B1(_i_CLEFIA128_state_reg _1), .O(n7784) );
  NR2GHD U11207 ( .I1(n7787), .I2(n7786), .O(n12303) );
  ND2HHD U11208 ( .I1(n13521), .I2(n7035), .O(n12086) );
  OAI12CHD U11209 ( .B1(n7035), .B2(n9807), .A1(n7254), .O(n7788) );
  NR2GHD U11210 ( .I1(n8533), .I2(n11706), .O(n8701) );
  XNR2HHD U11211 ( .I1(n13926), .I2(n13742), .O(n15520) );
  XNR2KHD U11212 ( .I1(n7790), .I2(n13925), .O(n14647) );
  XOR2HHD U11213 ( .I1(_i_CLEFIA128_keyL _76), .I2(n7792), .O(n7791) );
  ND3EHD U11214 ( .I1(n12832), .I2(n12790), .I3(n8232), .O(n7795) );
  OR2KHD U11215 ( .I1(n8315), .I2(n10206), .O(n8232) );
  ND2HHD U11216 ( .I1(n12674), .I2(n10905), .O(n7796) );
  OR2B1HHD U11217 ( .I1(n7216), .B1(n8199), .O(n10803) );
  XNR3EHD U11218 ( .I1(DOUT_66), .I2(n9978), .I3(n14993), .O(n10262) );
  AN2HHD U11219 ( .I1(n9249), .I2(n9242), .O(n9041) );
  OA12HHD U11220 ( .B1(n9122), .B2(n9120), .A1(n8264), .O(n7799) );
  ND2HHD U11221 ( .I1(n9980), .I2(n13608), .O(n7800) );
  OA13EHD U11222 ( .B1(n13140), .B2(n12026), .B3(n12025), .A1(n13622), .O(n7804) );
  AN2HHD U11223 ( .I1(n7805), .I2(n7004), .O(n11535) );
  ND2HHD U11224 ( .I1(n7807), .I2(n6982), .O(n13407) );
  AN2HHD U11225 ( .I1(n7807), .I2(n9343), .O(n13008) );
  NR2GHD U11226 ( .I1(n13006), .I2(n13007), .O(n7807) );
  BUFNHD U11227 ( .I(n9822), .O(n7808) );
  BUFNHD U11228 ( .I(n8992), .O(n7810) );
  ND2HHD U11229 ( .I1(n8583), .I2(n9621), .O(n8539) );
  ND2KHD U11230 ( .I1(n11681), .I2(n11794), .O(n9621) );
  XNR2KHD U11231 ( .I1(n7812), .I2(n11885), .O(n11904) );
  ND2HHD U11232 ( .I1(n11896), .I2(n7811), .O(n11903) );
  ND2KHD U11233 ( .I1(n7811), .I2(n11930), .O(n9214) );
  ND2HHD U11234 ( .I1(n9560), .I2(n6977), .O(n7814) );
  ND2HHD U11235 ( .I1(n12672), .I2(n6973), .O(n7815) );
  ND2HHD U11236 ( .I1(n7817), .I2(n10282), .O(n7816) );
  ND3EHD U11237 ( .I1(n7824), .I2(n12686), .I3(n7818), .O(n7817) );
  NR2GHD U11238 ( .I1(n12712), .I2(n9325), .O(n7821) );
  ND3EHD U11239 ( .I1(n12863), .I2(n7824), .I3(n7823), .O(n7822) );
  ND2KHD U11240 ( .I1(n10178), .I2(n9766), .O(n10798) );
  ND3EHD U11241 ( .I1(n12538), .I2(n10798), .I3(n12620), .O(n7826) );
  BUFNHD U11242 ( .I(n8164), .O(n7830) );
  NR2IHD U11243 ( .I1(n11893), .I2(n11911), .O(n8164) );
  ND2HHD U11244 ( .I1(n7831), .I2(n15500), .O(n15501) );
  ND2KHD U11245 ( .I1(n8797), .I2(_i_CLEFIA128_keyK _105), .O(n11879) );
  ND2HHD U11246 ( .I1(n9759), .I2(n7835), .O(n12161) );
  ND2KHD U11247 ( .I1(n9811), .I2(n9435), .O(n7835) );
  ND2DHD U11248 ( .I1(n7835), .I2(n13651), .O(n13830) );
  ND2CHD U11249 ( .I1(n7835), .I2(n8779), .O(n11724) );
  XOR2HHD U11250 ( .I1(n14332), .I2(n14331), .O(n7837) );
  ND2KHD U11251 ( .I1(n7041), .I2(n7808), .O(n9810) );
  ND2HHD U11252 ( .I1(n13829), .I2(n13652), .O(n9944) );
  ND2HHD U11253 ( .I1(n12066), .I2(n11713), .O(n13652) );
  ND3EHD U11254 ( .I1(n6985), .I2(n7020), .I3(n7843), .O(n12961) );
  NR3BHD U11255 ( .I1(n13809), .I2(n9525), .I3(n13807), .O(n7846) );
  OR2KHD U11256 ( .I1(n12238), .I2(n12237), .O(n8118) );
  ND2HHD U11257 ( .I1(n8887), .I2(n6635), .O(n7847) );
  AN2HHD U11258 ( .I1(n9335), .I2(n7848), .O(n9334) );
  ND2HHD U11259 ( .I1(n7219), .I2(_i_CLEFIA128_keyK _104), .O(n11869) );
  ND2HHD U11260 ( .I1(n9773), .I2(n12662), .O(n7849) );
  ND3EHD U11261 ( .I1(n8720), .I2(n8721), .I3(n11230), .O(n7850) );
  OAI12CHD U11262 ( .B1(n10808), .B2(n11203), .A1(n12646), .O(n7851) );
  ND2KHD U11263 ( .I1(n7854), .I2(n7852), .O(n8212) );
  ND3EHD U11264 ( .I1(n7855), .I2(n15247), .I3(_i_CLEFIA128_rndcnt_reg _0), .O(n10305) );
  AN3B1HHD U11265 ( .I1(n8789), .I2(n8198), .B1(n7866), .O(n10384) );
  ND3EHD U11266 ( .I1(n8035), .I2(n8032), .I3(n8496), .O(n7856) );
  ND2HHD U11267 ( .I1(n10319), .I2(_i_CLEFIA128_state_reg _1), .O(n7857) );
  ND2HHD U11268 ( .I1(n7859), .I2(n12312), .O(n9217) );
  AN2HHD U11269 ( .I1(n7860), .I2(n11201), .O(n8288) );
  NR2GHD U11270 ( .I1(n11061), .I2(n11060), .O(n7860) );
  ND2KHD U11271 ( .I1(n7254), .I2(n7809), .O(n13653) );
  AN2HHD U11272 ( .I1(n13506), .I2(n13550), .O(n8333) );
  ND2HHD U11273 ( .I1(n8832), .I2(n12296), .O(n7862) );
  ND2KHD U11274 ( .I1(n7386), .I2(n8209), .O(n12296) );
  ND2HHD U11275 ( .I1(n9811), .I2(n12145), .O(n8832) );
  ND2HHD U11276 ( .I1(n13646), .I2(n13653), .O(n13514) );
  OR2KHD U11277 ( .I1(n7863), .I2(n10332), .O(n7865) );
  ND3EHD U11278 ( .I1(n13138), .I2(n7867), .I3(n13601), .O(n13139) );
  ND3EHD U11279 ( .I1(n12943), .I2(n12942), .I3(n7867), .O(n12944) );
  XOR2HHD U11280 ( .I1(n10140), .I2(n6838), .O(n7868) );
  NR2GHD U11281 ( .I1(n12305), .I2(n8582), .O(n12316) );
  ND2KHD U11282 ( .I1(n13681), .I2(n12296), .O(n11804) );
  ND2HHD U11283 ( .I1(n7871), .I2(_i_CLEFIA128_state_reg _1), .O(n9720) );
  ND3EHD U11284 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(n11665), .I3(n15014), .O(n7871) );
  NR2IHD U11285 ( .I1(n7934), .I2(n11793), .O(n7933) );
  AN2HHD U11286 ( .I1(n11685), .I2(n10145), .O(n7872) );
  ND2KHD U11287 ( .I1(n9811), .I2(n7386), .O(n9612) );
  ND2HHD U11288 ( .I1(n9612), .I2(n13837), .O(n8834) );
  ND3EHD U11289 ( .I1(n9612), .I2(n9741), .I3(n13829), .O(n11708) );
  OA13EHD U11290 ( .B1(n7873), .B2(n11729), .B3(n11728), .A1(n13817), .O(n9829) );
  ND3EHD U11291 ( .I1(n9925), .I2(n11723), .I3(n10260), .O(n7873) );
  XOR2HHD U11292 ( .I1(n8762), .I2(n9923), .O(n14214) );
  ND2KHD U11293 ( .I1(n7291), .I2(n8204), .O(n7967) );
  ND2HHD U11294 ( .I1(n15392), .I2(n15380), .O(n15390) );
  XNR2KHD U11295 ( .I1(n13911), .I2(n13701), .O(n7985) );
  XOR2HHD U11296 ( .I1(n14243), .I2(n6816), .O(n13701) );
  XOR2HHD U11297 ( .I1(n14193), .I2(n9215), .O(n10116) );
  XNR2KHD U11298 ( .I1(n14106), .I2(n9519), .O(n9215) );
  XOR2HHD U11299 ( .I1(DOUT_68), .I2(n14332), .O(n10117) );
  ND2HHD U11300 ( .I1(n10561), .I2(n6560), .O(n7877) );
  NR2IHD U11301 ( .I1(n10431), .I2(n7879), .O(n10739) );
  INVCKGHD U11302 ( .I(n7884), .O(n7880) );
  ND3EHD U11303 ( .I1(n7881), .I2(n7883), .I3(n10968), .O(n8957) );
  AN3HHD U11304 ( .I1(n7884), .I2(n7885), .I3(n6975), .O(n7883) );
  ND2HHD U11305 ( .I1(n8888), .I2(n10959), .O(n7890) );
  ND2HHD U11306 ( .I1(n12448), .I2(n12479), .O(n7892) );
  ND2KHD U11307 ( .I1(n9903), .I2(n8768), .O(n12479) );
  ND2KHD U11308 ( .I1(n9087), .I2(n10599), .O(n12448) );
  ND2KHD U11309 ( .I1(n12484), .I2(n9800), .O(n9218) );
  ND2KHD U11310 ( .I1(n10978), .I2(n11439), .O(n11556) );
  ND2KHD U11311 ( .I1(n6873), .I2(n7671), .O(n11439) );
  ND2HHD U11312 ( .I1(n11554), .I2(n11555), .O(n7894) );
  ND2KHD U11313 ( .I1(n9903), .I2(n10599), .O(n11555) );
  ND2KHD U11314 ( .I1(n9194), .I2(n9903), .O(n11554) );
  ND2HHD U11315 ( .I1(n8797), .I2(_i_CLEFIA128_keyK _75), .O(n10418) );
  XOR2HHD U11316 ( .I1(n7896), .I2(n7985), .O(n8068) );
  XOR2HHD U11317 ( .I1(n14489), .I2(n8774), .O(n7896) );
  ND2KHD U11318 ( .I1(n7973), .I2(n7972), .O(n7977) );
  ND3EHD U11319 ( .I1(n7898), .I2(n10989), .I3(n7900), .O(n11311) );
  ND2HHD U11320 ( .I1(n7902), .I2(n7901), .O(n6187) );
  XNR2KHD U11321 ( .I1(n9215), .I2(n7903), .O(n10008) );
  XOR2HHD U11322 ( .I1(n14184), .I2(n9374), .O(n7903) );
  ND2HHD U11323 ( .I1(n8134), .I2(n8133), .O(n10205) );
  ND2HHD U11324 ( .I1(n8039), .I2(_i_CLEFIA128_keyK _83), .O(n9193) );
  AN2HHD U11325 ( .I1(n14043), .I2(n10296), .O(n8250) );
  AN2HHD U11326 ( .I1(n8227), .I2(n9455), .O(n7908) );
  OR3HHD U11327 ( .I1(n7912), .I2(n9953), .I3(n11177), .O(n11461) );
  ND2KHD U11328 ( .I1(n8237), .I2(n11417), .O(n9298) );
  ND2KHD U11329 ( .I1(n9017), .I2(n12484), .O(n11522) );
  ND3EHD U11330 ( .I1(n6961), .I2(n12297), .I3(n7918), .O(n7993) );
  ND2HHD U11331 ( .I1(n9650), .I2(n14076), .O(n7919) );
  ND2HHD U11332 ( .I1(n9551), .I2(n8329), .O(n7920) );
  ND3EHD U11333 ( .I1(n7923), .I2(n7922), .I3(DOUT_84), .O(n7924) );
  AN2HHD U11334 ( .I1(n13827), .I2(n7019), .O(n7925) );
  ND3EHD U11335 ( .I1(n8372), .I2(n9432), .I3(n6964), .O(n7928) );
  ND3EHD U11336 ( .I1(n12311), .I2(n12310), .I3(n13806), .O(n12314) );
  ND2HHD U11337 ( .I1(n7931), .I2(n8779), .O(n11716) );
  ND2HHD U11338 ( .I1(n7809), .I2(n7933), .O(n12088) );
  ND2HHD U11339 ( .I1(n7933), .I2(n12145), .O(n9309) );
  ND2HHD U11340 ( .I1(n7933), .I2(n8178), .O(n12150) );
  NR2GHD U11341 ( .I1(n7936), .I2(n8831), .O(n13827) );
  ND2HHD U11342 ( .I1(n6960), .I2(n9030), .O(n8831) );
  ND3EHD U11343 ( .I1(n13822), .I2(n8581), .I3(n13681), .O(n7936) );
  ND2HHD U11344 ( .I1(n12092), .I2(n13512), .O(n7938) );
  ND2HHD U11345 ( .I1(n7942), .I2(n13573), .O(n8605) );
  ND2DHD U11346 ( .I1(n7942), .I2(n7954), .O(n12101) );
  ND2CHD U11347 ( .I1(n7942), .I2(n12268), .O(n12036) );
  ND2CHD U11348 ( .I1(n7942), .I2(n12920), .O(n12281) );
  ND2CHD U11349 ( .I1(n7942), .I2(n13187), .O(n12271) );
  ND3CHD U11350 ( .I1(n12293), .I2(n9770), .I3(n7942), .O(n12294) );
  ND2KHD U11351 ( .I1(n13132), .I2(n10095), .O(n7942) );
  XOR2HHD U11352 ( .I1(n14994), .I2(n14351), .O(n14635) );
  XOR2HHD U11353 ( .I1(n13556), .I2(n14327), .O(n8830) );
  ND2KHD U11354 ( .I1(n14090), .I2(n7944), .O(n14351) );
  ND2HHD U11355 ( .I1(n7946), .I2(n7945), .O(n14994) );
  NR2GHD U11356 ( .I1(n13535), .I2(n13536), .O(n7946) );
  ND2HHD U11357 ( .I1(n7947), .I2(n13634), .O(n9879) );
  ND3EHD U11358 ( .I1(n7951), .I2(n7950), .I3(n7948), .O(n7947) );
  INVCKGHD U11359 ( .I(n12100), .O(n7949) );
  ND3EHD U11360 ( .I1(n12928), .I2(n13211), .I3(n12109), .O(n13631) );
  ND2HHD U11361 ( .I1(n7953), .I2(n8262), .O(n6274) );
  ND2HHD U11362 ( .I1(n7952), .I2(n7043), .O(n7953) );
  XOR2HHD U11363 ( .I1(n12138), .I2(n10000), .O(n9540) );
  AN2HHD U11364 ( .I1(n7954), .I2(n13577), .O(n8443) );
  ND2CHD U11365 ( .I1(n7954), .I2(n13125), .O(n12059) );
  ND2CHD U11366 ( .I1(n7954), .I2(n13592), .O(n13171) );
  ND2KHD U11367 ( .I1(n11997), .I2(n12915), .O(n7954) );
  BUFMHD U11368 ( .I(n13556), .O(n7955) );
  ND2HHD U11369 ( .I1(n8729), .I2(n13208), .O(n12921) );
  NR2GHD U11370 ( .I1(n10006), .I2(n7962), .O(n7961) );
  ND3EHD U11371 ( .I1(n6835), .I2(n13211), .I3(n7964), .O(n7962) );
  OR2CHD U11372 ( .I1(n12377), .I2(n8881), .O(n7964) );
  ND2HHD U11373 ( .I1(n8597), .I2(n7966), .O(n8596) );
  ND3EHD U11374 ( .I1(n9576), .I2(n7966), .I3(n9578), .O(n13245) );
  AN2HHD U11375 ( .I1(n12127), .I2(n7968), .O(n13184) );
  XNR3EHD U11376 ( .I1(n7971), .I2(n13267), .I3(n9893), .O(n7998) );
  XOR2HHD U11377 ( .I1(n8719), .I2(n9637), .O(n9893) );
  XOR2HHD U11378 ( .I1(n9959), .I2(n9914), .O(n13267) );
  XNR3EHD U11379 ( .I1(DOUT_19), .I2(n14167), .I3(n9896), .O(n7971) );
  ND3EHD U11380 ( .I1(n6925), .I2(n7389), .I3(n11592), .O(n7976) );
  ND2HHD U11381 ( .I1(n7974), .I2(n7976), .O(n7975) );
  OR3HHD U11382 ( .I1(n10948), .I2(n7981), .I3(n10821), .O(n7980) );
  ND2HHD U11383 ( .I1(n7982), .I2(n10960), .O(n7981) );
  ND3EHD U11384 ( .I1(n7983), .I2(n15140), .I3(_i_CLEFIA128_rndcnt_reg _0), .O(n11589) );
  XOR2HHD U11385 ( .I1(n6725), .I2(n8549), .O(n15269) );
  ND2HHD U11386 ( .I1(n7986), .I2(n11523), .O(n11153) );
  NR2GHD U11387 ( .I1(n9900), .I2(n9901), .O(n7986) );
  INVGHD U11388 ( .I(n7988), .O(n7987) );
  NR2IHD U11389 ( .I1(n9941), .I2(n11662), .O(n7988) );
  ND2CHD U11390 ( .I1(n7990), .I2(n8237), .O(n10615) );
  ND2KHD U11391 ( .I1(n8899), .I2(n8379), .O(n8577) );
  OR2KHD U11392 ( .I1(n6832), .I2(n12748), .O(n7991) );
  OR3HHD U11393 ( .I1(n13836), .I2(n9835), .I3(n9944), .O(n12168) );
  ND3EHD U11394 ( .I1(n12149), .I2(n8252), .I3(n13818), .O(n7996) );
  ND3EHD U11395 ( .I1(n12148), .I2(n12321), .I3(n10142), .O(n7997) );
  XNR2KHD U11396 ( .I1(n14367), .I2(n14366), .O(n9895) );
  ND2HHD U11397 ( .I1(n7999), .I2(n8000), .O(n6177) );
  ND2HHD U11398 ( .I1(n10465), .I2(n7389), .O(n10243) );
  INVCKGHD U11399 ( .I(n11332), .O(n8002) );
  ND2HHD U11400 ( .I1(n8484), .I2(n11376), .O(n8003) );
  NR2GHD U11401 ( .I1(n8004), .I2(n8005), .O(n8484) );
  ND2HHD U11402 ( .I1(n11098), .I2(n11097), .O(n8005) );
  ND2DHD U11403 ( .I1(n6887), .I2(n7043), .O(n8007) );
  ND3EHD U11404 ( .I1(n8008), .I2(n8010), .I3(n15320), .O(n6116) );
  ND2HHD U11405 ( .I1(n8009), .I2(n15321), .O(n8008) );
  NR2GHD U11406 ( .I1(n6951), .I2(n8013), .O(n11015) );
  ND2KHD U11407 ( .I1(n8176), .I2(n7548), .O(n8012) );
  ND2HHD U11408 ( .I1(n6947), .I2(n11508), .O(n8016) );
  ND2HHD U11409 ( .I1(n8247), .I2(n6944), .O(n8017) );
  OA13EHD U11410 ( .B1(n12557), .B2(n11517), .B3(n12592), .A1(n12575), .O(n11518) );
  NR2IHD U11411 ( .I1(_i_CLEFIA128_keyK _67), .I2(n15304), .O(n8021) );
  NR2GHD U11412 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(n8021), .O(n8020) );
  ND2KHD U11413 ( .I1(n8023), .I2(n8022), .O(n10198) );
  AN2HHD U11414 ( .I1(n8028), .I2(n8025), .O(n13072) );
  ND2HHD U11415 ( .I1(n11834), .I2(n8027), .O(n8026) );
  ND2KHD U11416 ( .I1(n9597), .I2(n8078), .O(n13053) );
  NR2GHD U11417 ( .I1(n9920), .I2(n12195), .O(n8028) );
  ND2KHD U11418 ( .I1(n11818), .I2(n6837), .O(n9631) );
  ND2HHD U11419 ( .I1(n9074), .I2(n9073), .O(n8756) );
  ND2HHD U11420 ( .I1(n8899), .I2(n8345), .O(n8033) );
  XNR2KHD U11421 ( .I1(n8037), .I2(n8036), .O(n15503) );
  XOR2HHD U11422 ( .I1(n13912), .I2(n14804), .O(n8037) );
  ND3EHD U11423 ( .I1(n8038), .I2(n14953), .I3(_i_CLEFIA128_rndcnt_reg _0), .O(n10323) );
  ND2HHD U11424 ( .I1(n8041), .I2(n8040), .O(n11057) );
  ND2KHD U11425 ( .I1(n6842), .I2(n6883), .O(n12652) );
  ND2KHD U11426 ( .I1(n9680), .I2(n10874), .O(n11250) );
  ND3EHD U11427 ( .I1(n8045), .I2(n8044), .I3(_i_CLEFIA128_rndcnt_reg _0), .O(n8047) );
  ND2HHD U11428 ( .I1(_i_CLEFIA128_keyL _61), .I2(n9494), .O(n8044) );
  ND3EHD U11429 ( .I1(n11564), .I2(n8047), .I3(_i_CLEFIA128_state_reg _1), .O(n11565) );
  INVKHD U11430 ( .I(n8048), .O(n8198) );
  ND2HHD U11431 ( .I1(n8050), .I2(n6996), .O(n8049) );
  ND2HHD U11432 ( .I1(n10286), .I2(n9683), .O(n8050) );
  NR2IHD U11433 ( .I1(n8798), .I2(n8051), .O(n8052) );
  INVQHD U11434 ( .I(_i_CLEFIA128_keyK _89), .O(n8051) );
  XNR2HHD U11435 ( .I1(_i_CLEFIA128_keyL _89), .I2(n8052), .O(n9950) );
  OR2EHD U11436 ( .I1(n10002), .I2(n12184), .O(n8054) );
  OA13EHD U11437 ( .B1(n8056), .B2(n8057), .B3(n12188), .A1(n14087), .O(n8055));
  OA13EHD U11438 ( .B1(n12212), .B2(n12213), .B3(n8059), .A1(n14067), .O(n8058) );
  ND2CHD U11439 ( .I1(n6587), .I2(n7842), .O(n12194) );
  ND2KHD U11440 ( .I1(n8204), .I2(n8078), .O(n8061) );
  XOR2HHD U11441 ( .I1(n10127), .I2(n8062), .O(n9697) );
  XOR2HHD U11442 ( .I1(n14184), .I2(n8063), .O(n8062) );
  OR3HHD U11443 ( .I1(n11630), .I2(n8997), .I3(n13080), .O(n12185) );
  ND2HHD U11444 ( .I1(n13096), .I2(n13469), .O(n8073) );
  INVCKGHD U11445 ( .I(n13075), .O(n8069) );
  ND2HHD U11446 ( .I1(n15067), .I2(n15500), .O(n8075) );
  ND2HHD U11447 ( .I1(n9994), .I2(n8827), .O(n8077) );
  ND2KHD U11448 ( .I1(n8204), .I2(n6837), .O(n8190) );
  NR2GHD U11449 ( .I1(n8080), .I2(n11745), .O(n13062) );
  ND3EHD U11450 ( .I1(n8190), .I2(n11744), .I3(n12208), .O(n8080) );
  ND2HHD U11451 ( .I1(n7034), .I2(n8078), .O(n11744) );
  NR2IHD U11452 ( .I1(n8798), .I2(n8081), .O(n8082) );
  XOR2HHD U11453 ( .I1(_i_CLEFIA128_keyL _121), .I2(n8082), .O(n9995) );
  ND2KHD U11454 ( .I1(n11707), .I2(n11679), .O(n8083) );
  ND2HHD U11455 ( .I1(n12321), .I2(n13818), .O(n8085) );
  NR2GHD U11456 ( .I1(n6785), .I2(n8195), .O(n12152) );
  ND2HHD U11457 ( .I1(n8628), .I2(n13671), .O(n12151) );
  NR2GHD U11458 ( .I1(n12317), .I2(n12318), .O(n8086) );
  ND2HHD U11459 ( .I1(n13652), .I2(n13842), .O(n12317) );
  ND2HHD U11460 ( .I1(n9621), .I2(n13821), .O(n12318) );
  ND3EHD U11461 ( .I1(n8090), .I2(n14114), .I3(n8087), .O(n6171) );
  ND2HHD U11462 ( .I1(n15095), .I2(n11130), .O(n8087) );
  XNR3EHD U11463 ( .I1(n14109), .I2(n14108), .I3(n14107), .O(n8088) );
  XNR2KHD U11464 ( .I1(n8092), .I2(n8091), .O(n15235) );
  XNR2HHD U11465 ( .I1(n14803), .I2(n14804), .O(n8092) );
  ND2HHD U11466 ( .I1(n11834), .I2(n9628), .O(n13217) );
  INVCHD U11467 ( .I(n8094), .O(n11164) );
  ND2HHD U11468 ( .I1(n6999), .I2(n8093), .O(n10723) );
  ND2HHD U11469 ( .I1(n8797), .I2(_i_CLEFIA128_keyK _17), .O(n8099) );
  ND2HHD U11470 ( .I1(n8097), .I2(_i_CLEFIA128_state_reg _1), .O(n8096) );
  ND2HHD U11471 ( .I1(n8101), .I2(n11482), .O(n11483) );
  ND3EHD U11472 ( .I1(n12582), .I2(n12737), .I3(n8101), .O(n9417) );
  ND3EHD U11473 ( .I1(n12749), .I2(n8101), .I3(n12765), .O(n12720) );
  ND2KHD U11474 ( .I1(n8182), .I2(n9738), .O(n8101) );
  OR3HHD U11475 ( .I1(_i_CLEFIA128_keyL _0), .I2(n8102), .I3(n8589), .O(n8103) );
  ND2HHD U11476 ( .I1(n8797), .I2(_i_CLEFIA128_rndcnt_reg _0), .O(n8105) );
  ND2HHD U11477 ( .I1(_i_CLEFIA128_keyK _0), .I2(_i_CLEFIA128_keyL _0), .O(n8106) );
  INVCKGHD U11478 ( .I(n8108), .O(n8107) );
  NR2GHD U11479 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(n8111), .O(n8110) );
  NR2IHD U11480 ( .I1(n10209), .I2(n8114), .O(n11895) );
  NR2BHD U11481 ( .I1(n12328), .I2(n8114), .O(n12330) );
  ND2HHD U11482 ( .I1(n11852), .I2(n7842), .O(n9315) );
  AN3HHD U11483 ( .I1(n10225), .I2(n9568), .I3(n7977), .O(n8227) );
  ND2HHD U11484 ( .I1(n8515), .I2(n8018), .O(n8117) );
  NR2IHD U11485 ( .I1(n7674), .I2(n11504), .O(n12562) );
  NR2IHD U11486 ( .I1(n8798), .I2(n8121), .O(n8122) );
  INVQHD U11487 ( .I(_i_CLEFIA128_keyK _114), .O(n8121) );
  ND2HHD U11488 ( .I1(n9125), .I2(n8123), .O(n9274) );
  ND2HHD U11489 ( .I1(n11863), .I2(n11861), .O(n8125) );
  ND2HHD U11490 ( .I1(n8845), .I2(n8126), .O(n8833) );
  AN2KHD U11491 ( .I1(n11640), .I2(n13216), .O(n14076) );
  ND3EHD U11492 ( .I1(n11820), .I2(n14080), .I3(n8197), .O(n8129) );
  ND2KHD U11493 ( .I1(n9628), .I2(n6837), .O(n8197) );
  OA12HHD U11494 ( .B1(n11595), .B2(_i_CLEFIA128_keyL _127), .A1(n6927), .O(n8131) );
  OR2KHD U11495 ( .I1(n10446), .I2(n8133), .O(n10761) );
  ND2KHD U11496 ( .I1(n12291), .I2(n8185), .O(n13614) );
  ND2HHD U11497 ( .I1(n12291), .I2(n12383), .O(n13582) );
  ND2KHD U11498 ( .I1(n10169), .I2(n10168), .O(n8136) );
  ND2KHD U11499 ( .I1(n8136), .I2(n10659), .O(n10328) );
  OR2CHD U11500 ( .I1(n11260), .I2(n12658), .O(n10681) );
  ND2HHD U11501 ( .I1(n8138), .I2(n10171), .O(n10170) );
  ND2KHD U11502 ( .I1(n10855), .I2(n10847), .O(n11260) );
  ND2KHD U11503 ( .I1(n11175), .I2(n7040), .O(n11548) );
  ND2HHD U11504 ( .I1(n8140), .I2(n8303), .O(n12716) );
  NR2GHD U11505 ( .I1(n8139), .I2(n7030), .O(n8303) );
  ND2HHD U11506 ( .I1(n12674), .I2(n8812), .O(n8139) );
  ND3EHD U11507 ( .I1(n8141), .I2(n8146), .I3(n8144), .O(n12667) );
  NR2GHD U11508 ( .I1(n8143), .I2(n8142), .O(n8141) );
  ND2HHD U11509 ( .I1(n9735), .I2(n10888), .O(n8143) );
  INVCKGHD U11510 ( .I(n12799), .O(n8146) );
  ND3EHD U11511 ( .I1(n8149), .I2(n8316), .I3(n8147), .O(n11824) );
  OR3HHD U11512 ( .I1(n11819), .I2(n8148), .I3(n13232), .O(n14084) );
  ND2HHD U11513 ( .I1(n9006), .I2(n11820), .O(n8150) );
  OAI112BHD U11514 ( .C1(n11603), .C2(n15233), .A1(n11608), .B1(n8152), .O(n8151) );
  ND3EHD U11515 ( .I1(n8158), .I2(n8157), .I3(n8156), .O(n8154) );
  ND3EHD U11516 ( .I1(n8162), .I2(n8160), .I3(n8689), .O(n8155) );
  AN2HHD U11517 ( .I1(n10113), .I2(n11989), .O(n8161) );
  ND2HHD U11518 ( .I1(n8692), .I2(n10112), .O(n8162) );
  ND2HHD U11519 ( .I1(n8163), .I2(n14255), .O(n6122) );
  OA12HHD U11520 ( .B1(n9895), .B2(n15513), .A1(n15489), .O(n8168) );
  ND2HHD U11521 ( .I1(n9272), .I2(n9273), .O(n8170) );
  ND2HHD U11522 ( .I1(n8171), .I2(n9906), .O(n9905) );
  ND3EHD U11523 ( .I1(n9275), .I2(n9276), .I3(n9907), .O(n8171) );
  ND2HHD U11524 ( .I1(n8172), .I2(n7389), .O(n9907) );
  XOR2HHD U11525 ( .I1(_i_CLEFIA128_keyL _85), .I2(n10556), .O(n8172) );
  AN3HHD U11526 ( .I1(n9667), .I2(n8383), .I3(n14063), .O(n11770) );
  AN2HHD U11527 ( .I1(n11744), .I2(n14072), .O(n8383) );
  AN2EHD U11528 ( .I1(n12120), .I2(n9456), .O(n8223) );
  XOR2HHD U11529 ( .I1(n14329), .I2(n9978), .O(n12445) );
  ND3HHD U11530 ( .I1(n11253), .I2(n10847), .I3(n11233), .O(n10647) );
  ND2HHD U11531 ( .I1(n9096), .I2(n13426), .O(n10101) );
  NR2IHD U11532 ( .I1(n9824), .I2(n9829), .O(n9803) );
  AN2EHD U11533 ( .I1(n9207), .I2(n12120), .O(n8228) );
  ND2KHD U11534 ( .I1(n8798), .I2(_i_CLEFIA128_keyL _64), .O(n9014) );
  NR2GHD U11535 ( .I1(n13689), .I2(n13688), .O(n13690) );
  ND2KHD U11536 ( .I1(n12181), .I2(n11820), .O(n13235) );
  ND2KHD U11537 ( .I1(n9183), .I2(n7034), .O(n12181) );
  ND2KHD U11538 ( .I1(n7907), .I2(n8204), .O(n11820) );
  OR3EHD U11539 ( .I1(n12525), .I2(n12524), .I3(n12523), .O(n12527) );
  ND3HHD U11540 ( .I1(n13589), .I2(n6897), .I3(n8657), .O(n13165) );
  ND2HHD U11541 ( .I1(n8116), .I2(n9898), .O(n8483) );
  ND2HHD U11542 ( .I1(n12562), .I2(n9049), .O(n8470) );
  ND2KHD U11543 ( .I1(n9587), .I2(n12431), .O(n12224) );
  AN2HHD U11544 ( .I1(n13440), .I2(n13444), .O(n13389) );
  ND2DHD U11545 ( .I1(n9102), .I2(n8697), .O(n8696) );
  ND2KHD U11546 ( .I1(n9831), .I2(n9606), .O(n8757) );
  INVQHD U11547 ( .I(_i_CLEFIA128_keyL _5), .O(n15257) );
  ND2HHD U11548 ( .I1(n8637), .I2(n12671), .O(n8636) );
  ND2KHD U11549 ( .I1(n13521), .I2(n7810), .O(n12163) );
  AN3HHD U11550 ( .I1(n10960), .I2(n6734), .I3(n12868), .O(n10890) );
  ND2KHD U11551 ( .I1(n10746), .I2(n8215), .O(n12868) );
  OR3HHD U11552 ( .I1(n12703), .I2(n12701), .I3(n12702), .O(n12707) );
  ND2DHD U11553 ( .I1(n12714), .I2(n7033), .O(n12702) );
  NR2EHD U11554 ( .I1(n12809), .I2(n8427), .O(n12788) );
  ND2KHD U11555 ( .I1(n8191), .I2(n7723), .O(n8547) );
  ND2KHD U11556 ( .I1(n11995), .I2(n8185), .O(n9998) );
  ND2HHD U11557 ( .I1(n8572), .I2(n7389), .O(n8556) );
  INVQHD U11558 ( .I(n8854), .O(n10794) );
  ND2DHD U11559 ( .I1(n9832), .I2(n13572), .O(n10224) );
  NR2GHD U11560 ( .I1(n11722), .I2(n9926), .O(n9925) );
  NR2EHD U11561 ( .I1(n12330), .I2(n12329), .O(n13397) );
  BUFQHD U11562 ( .I(n11898), .O(n12226) );
  ND2HHD U11563 ( .I1(n9605), .I2(n14070), .O(n13488) );
  OA12EHD U11564 ( .B1(n14647), .B2(n15512), .A1(n14646), .O(n14648) );
  AN3HHD U11565 ( .I1(n8470), .I2(n12731), .I3(n11511), .O(n12740) );
  ND2KHD U11566 ( .I1(n9099), .I2(n6832), .O(n10474) );
  ND2KHD U11567 ( .I1(n8200), .I2(n8196), .O(n12320) );
  ND3EHD U11568 ( .I1(n12543), .I2(n12542), .I3(n12541), .O(n12544) );
  NR2IHD U11569 ( .I1(n9668), .I2(n11490), .O(n9074) );
  NR2GHD U11570 ( .I1(n12314), .I2(n9032), .O(n8894) );
  ND3EHD U11571 ( .I1(n12832), .I2(n12674), .I3(n12673), .O(n8926) );
  OR3EHD U11572 ( .I1(n10677), .I2(n12510), .I3(n10678), .O(n10685) );
  NR2GHD U11573 ( .I1(n13473), .I2(n8595), .O(n8643) );
  ND2HHD U11574 ( .I1(n12241), .I2(n9620), .O(n13427) );
  ND3EHD U11575 ( .I1(n9345), .I2(n12814), .I3(n10283), .O(n8637) );
  ND2HHD U11576 ( .I1(n8583), .I2(n13821), .O(n12307) );
  ND2KHD U11577 ( .I1(n10219), .I2(n8215), .O(n8495) );
  ND2KHD U11578 ( .I1(n8618), .I2(n8617), .O(n8624) );
  NR2IHD U11579 ( .I1(n8693), .I2(n11706), .O(n8618) );
  ND2HHD U11580 ( .I1(n8916), .I2(n10741), .O(n12673) );
  OA112HHD U11581 ( .C1(n9414), .C2(n10032), .A1(n9413), .B1(n10028), .O(n10326) );
  ND2KHD U11582 ( .I1(n7034), .I2(n6837), .O(n11646) );
  NR2IHD U11583 ( .I1(n7897), .I2(n11762), .O(n12190) );
  OA12EHD U11584 ( .B1(n15336), .B2(n15335), .A1(n15333), .O(n8855) );
  BUFMHD U11585 ( .I(n10419), .O(n10442) );
  ND2HHD U11586 ( .I1(n9074), .I2(n9073), .O(n14243) );
  ND2DHD U11587 ( .I1(n6694), .I2(n12092), .O(n8846) );
  ND2KHD U11588 ( .I1(n9811), .I2(n7809), .O(n12092) );
  BUFQHD U11589 ( .I(n9961), .O(n8179) );
  BUFQHD U11590 ( .I(n11090), .O(n8180) );
  ND3EHD U11591 ( .I1(n13969), .I2(n13968), .I3(n13967), .O(n6173) );
  ND2HHD U11592 ( .I1(n15367), .I2(n11130), .O(n13967) );
  NR2GHD U11593 ( .I1(n9188), .I2(n8990), .O(n9165) );
  INVNHD U11594 ( .I(n9188), .O(n9580) );
  ND2KHD U11595 ( .I1(n6881), .I2(n9189), .O(n9188) );
  INVQHD U11596 ( .I(n8184), .O(n8185) );
  ND2HHD U11597 ( .I1(n8285), .I2(n9316), .O(n13095) );
  ND2KHD U11598 ( .I1(n9841), .I2(n10259), .O(n12748) );
  ND2HHD U11599 ( .I1(n11772), .I2(n14087), .O(n9228) );
  BUFQHD U11600 ( .I(n10334), .O(n8189) );
  NR2IHD U11601 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(n8797), .O(n10334) );
  BUFQHD U11602 ( .I(n8991), .O(n8191) );
  INVMHD U11603 ( .I(_i_CLEFIA128_keyL _72), .O(n15189) );
  ND2DHD U11604 ( .I1(n15235), .I2(n11130), .O(n14112) );
  ND2KHD U11605 ( .I1(n11634), .I2(n11614), .O(n12189) );
  INVQHD U11606 ( .I(n8195), .O(n8196) );
  ND2KHD U11607 ( .I1(n9581), .I2(n8191), .O(n8977) );
  XNR2HHD U11608 ( .I1(n14634), .I2(n14635), .O(n9743) );
  INVNHD U11609 ( .I(n8203), .O(n8204) );
  INVDHD U11610 ( .I(n14246), .O(n9870) );
  INVJHD U11611 ( .I(n12952), .O(n12346) );
  ND3CHD U11612 ( .I1(n8973), .I2(n7389), .I3(n8975), .O(n8972) );
  XNR2HHD U11613 ( .I1(_i_CLEFIA128_CON_T_xi _11), .I2(DOUT_36), .O(n9442));
  INVDHD U11614 ( .I(n10469), .O(n10071) );
  NR2GHD U11615 ( .I1(n10051), .I2(n11811), .O(n12066) );
  MUX2CHD U11616 ( .A(n10401), .B(n10400), .S(_i_CLEFIA128_keyL _79), .O(n10406) );
  NR2BHD U11617 ( .I1(n10399), .I2(n8189), .O(n10401) );
  ND2CHD U11618 ( .I1(n8224), .I2(_i_CLEFIA128_keyK _79), .O(n10400) );
  NR2CHD U11619 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(_i_CLEFIA128_keyK _79), .O(n10399) );
  ND2HHD U11620 ( .I1(n7808), .I2(n9549), .O(n11678) );
  ND2DHD U11621 ( .I1(n12012), .I2(n9478), .O(n9477) );
  MUX2CHD U11622 ( .A(n12009), .B(n12008), .S(_i_CLEFIA128_keyL _103), .O(n12013) );
  INVDHD U11623 ( .I(n6734), .O(n8970) );
  NR2GHD U11624 ( .I1(n10666), .I2(n10665), .O(n12546) );
  ND3CHD U11625 ( .I1(n11419), .I2(n7900), .I3(n9222), .O(n11421) );
  ND2HHD U11626 ( .I1(n12393), .I2(n13590), .O(n12117) );
  INVKHD U11627 ( .I(n9015), .O(n13175) );
  ND2CHD U11628 ( .I1(n13121), .I2(n13614), .O(n12262) );
  NR2CHD U11629 ( .I1(n9173), .I2(n14444), .O(n10299) );
  ND2HHD U11630 ( .I1(n9270), .I2(_i_CLEFIA128_state_reg _0), .O(n14719) );
  OA22CHD U11631 ( .A1(n15344), .A2(n15420), .B1(n15352), .B2(n13288), .O(n14537) );
  OA22CHD U11632 ( .A1(n9528), .A2(n15420), .B1(n15029), .B2(n13339), .O(n14638) );
  OA22CHD U11633 ( .A1(n15258), .A2(n15416), .B1(n13339), .B2(n15281), .O(n15259) );
  OA22CHD U11634 ( .A1(n15360), .A2(n15416), .B1(n13339), .B2(n15274), .O(n14858) );
  OA22CHD U11635 ( .A1(n15316), .A2(n15416), .B1(n13339), .B2(n15179), .O(n15180) );
  OA22CHD U11636 ( .A1(n15185), .A2(n15420), .B1(n15189), .B2(n13339), .O(n14897) );
  OA22CHD U11637 ( .A1(n15475), .A2(n15416), .B1(n13339), .B2(n7143), .O(n14824) );
  OA22CHD U11638 ( .A1(n14828), .A2(n15416), .B1(n13339), .B2(n14936), .O(n14829) );
  OA22CHD U11639 ( .A1(n14871), .A2(n15416), .B1(n13339), .B2(n15403), .O(n14872) );
  OA22CHD U11640 ( .A1(n15300), .A2(n15420), .B1(n14988), .B2(n13339), .O(n14990) );
  OA22CHD U11641 ( .A1(n15304), .A2(n15420), .B1(n14991), .B2(n13339), .O(n14592) );
  OA22CHD U11642 ( .A1(n15223), .A2(n15416), .B1(n13339), .B2(n15306), .O(n14968) );
  OA22CHD U11643 ( .A1(n15442), .A2(n15416), .B1(n13339), .B2(n15073), .O(n14973) );
  INVCHD U11644 ( .I(n14444), .O(n14403) );
  OR2CHD U11645 ( .I1(n15124), .I2(n15422), .O(n15118) );
  OA112CHD U11646 ( .C1(n15420), .C2(n15243), .A1(n15117), .B1(n15116), .O(n15119) );
  ND2CHD U11647 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _84), .O(n15117) );
  OR2CHD U11648 ( .I1(n15290), .I2(n15422), .O(n15291) );
  ND2CHD U11649 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _69), .O(n15288) );
  OR2CHD U11650 ( .I1(n14954), .I2(n15422), .O(n14955) );
  OA112CHD U11651 ( .C1(n15420), .C2(n14953), .A1(n14952), .B1(n14951), .O(n14956) );
  ND2CHD U11652 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _89), .O(n14952) );
  OA112CHD U11653 ( .C1(n14742), .C2(n14469), .A1(n14718), .B1(n14447), .O(n14448) );
  ND2CHD U11654 ( .I1(n14446), .I2(_i_CLEFIA128_CON_T_x _0), .O(n14447) );
  ND2CHD U11655 ( .I1(n14432), .I2(n14445), .O(n14446) );
  XOR2HHD U11656 ( .I1(_i_CLEFIA128_keyL _120), .I2(n11591), .O(n11592) );
  ND2DHD U11657 ( .I1(n8973), .I2(n7389), .O(n8941) );
  ND2HHD U11658 ( .I1(n9274), .I2(n9269), .O(n9267) );
  NR2EHD U11659 ( .I1(n9270), .I2(n11864), .O(n9269) );
  INVDHD U11660 ( .I(n10411), .O(n9447) );
  ND2DHD U11661 ( .I1(n6878), .I2(n6796), .O(n9323) );
  ND2DHD U11662 ( .I1(n13096), .I2(n13469), .O(n8649) );
  ND3CHD U11663 ( .I1(n11881), .I2(_i_CLEFIA128_rndcnt_reg _0), .I3(n15124), .O(n11882) );
  OR2EHD U11664 ( .I1(n14707), .I2(n8680), .O(n8429) );
  ND2HHD U11665 ( .I1(n12427), .I2(n13372), .O(n9937) );
  ND3CHD U11666 ( .I1(n13652), .I2(n12159), .I3(n11806), .O(n11807) );
  NR2EHD U11667 ( .I1(n8841), .I2(n12161), .O(n8840) );
  ND2DHD U11668 ( .I1(n13088), .I2(n13098), .O(n13067) );
  ND2HHD U11669 ( .I1(n9342), .I2(n13004), .O(n9387) );
  INVKHD U11670 ( .I(n9256), .O(n10712) );
  ND2DHD U11671 ( .I1(n6883), .I2(n12638), .O(n12518) );
  AN2HHD U11672 ( .I1(n10893), .I2(n12796), .O(n8921) );
  ND2CHD U11673 ( .I1(n7723), .I2(n12794), .O(n10962) );
  NR2GHD U11674 ( .I1(n9488), .I2(n9489), .O(n13106) );
  ND2HHD U11675 ( .I1(n9462), .I2(n9806), .O(n8595) );
  ND2HHD U11676 ( .I1(n9694), .I2(n8188), .O(n11323) );
  NR2BHD U11677 ( .I1(n10335), .I2(n8189), .O(n10336) );
  NR2CHD U11678 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(_i_CLEFIA128_keyK _94), .O(n10335) );
  ND2CHD U11679 ( .I1(n11505), .I2(n6833), .O(n10472) );
  NR2BHD U11680 ( .I1(n12117), .I2(n12039), .O(n12040) );
  NR2BHD U11681 ( .I1(n11594), .I2(n8189), .O(n11595) );
  NR2CHD U11682 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(_i_CLEFIA128_keyK _127), .O(n11594) );
  ND2DHD U11683 ( .I1(n12559), .I2(n12765), .O(n11017) );
  NR2CHD U11684 ( .I1(n12757), .I2(n11033), .O(n11037) );
  ND2HHD U11685 ( .I1(n9300), .I2(n12302), .O(n9299) );
  ND2CHD U11686 ( .I1(n11403), .I2(n12586), .O(n11350) );
  ND3CHD U11687 ( .I1(n12621), .I2(n12521), .I3(n12635), .O(n10649) );
  AN3EHD U11688 ( .I1(n13024), .I2(n13447), .I3(n12350), .O(n12247) );
  ND2DHD U11689 ( .I1(n9152), .I2(n12089), .O(n11784) );
  ND3CHD U11690 ( .I1(n9806), .I2(n14043), .I3(n13222), .O(n11826) );
  INVDHD U11691 ( .I(n12935), .O(n8892) );
  ND2HHD U11692 ( .I1(n13194), .I2(n6897), .O(n12104) );
  NR2EHD U11693 ( .I1(n12744), .I2(n12745), .O(n8684) );
  ND2HHD U11694 ( .I1(n12722), .I2(n12719), .O(n8460) );
  ND2DHD U11695 ( .I1(n12479), .I2(n11459), .O(n9900) );
  ND2DHD U11696 ( .I1(n11155), .I2(n9298), .O(n11158) );
  NR2CHD U11697 ( .I1(n10026), .I2(n13836), .O(n8736) );
  ND2DHD U11698 ( .I1(n9604), .I2(n9435), .O(n12080) );
  ND2CHD U11699 ( .I1(n12163), .I2(n12069), .O(n12071) );
  ND2CHD U11700 ( .I1(n13506), .I2(n13829), .O(n12070) );
  NR2EHD U11701 ( .I1(n9259), .I2(n6726), .O(n9258) );
  ND2DHD U11702 ( .I1(n8962), .I2(n8977), .O(n10729) );
  ND3CHD U11703 ( .I1(n8391), .I2(n9886), .I3(n13125), .O(n12396) );
  NR2EHD U11704 ( .I1(n12404), .I2(n12921), .O(n12259) );
  ND2DHD U11705 ( .I1(n13125), .I2(n9639), .O(n12256) );
  ND2CHD U11706 ( .I1(n12619), .I2(n12609), .O(n11249) );
  NR2BHD U11707 ( .I1(n10344), .I2(n8189), .O(n10346) );
  NR2CHD U11708 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(_i_CLEFIA128_keyK _95), .O(n10344) );
  ND3CHD U11709 ( .I1(n8376), .I2(n13589), .I3(n8866), .O(n12058) );
  OA13EHD U11710 ( .B1(n10718), .B2(n11467), .B3(n10985), .A1(n12462), .O(n10727) );
  ND3CHD U11711 ( .I1(n13167), .I2(n8715), .I3(n13168), .O(n8714) );
  INVDHD U11712 ( .I(n8786), .O(n8746) );
  NR2GHD U11713 ( .I1(n11389), .I2(n11390), .O(n10089) );
  OA22CHD U11714 ( .A1(n15373), .A2(n15416), .B1(n13339), .B2(n15121), .O(n15122) );
  OA22CHD U11715 ( .A1(n15115), .A2(n15416), .B1(n13339), .B2(n15125), .O(n15116) );
  ND2CHD U11716 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _105), .O(n14602) );
  OA22CHD U11717 ( .A1(n15242), .A2(n15420), .B1(n15247), .B2(n13339), .O(n14603) );
  ND2CHD U11718 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _112), .O(n15230) );
  ND2CHD U11719 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _119), .O(n15097) );
  OA22CHD U11720 ( .A1(n15494), .A2(n15416), .B1(n13339), .B2(n15233), .O(n15085) );
  OA22CHD U11721 ( .A1(n15432), .A2(n15416), .B1(n13339), .B2(n15100), .O(n13340) );
  ND2CHD U11722 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _126), .O(n14510) );
  OA22CHD U11723 ( .A1(n15092), .A2(n15420), .B1(n13339), .B2(n9474), .O(n14511) );
  OA22CHD U11724 ( .A1(n15498), .A2(n15416), .B1(n13339), .B2(n15239), .O(n15081) );
  OA22CHD U11725 ( .A1(n15437), .A2(n15416), .B1(n13339), .B2(n15249), .O(n15102) );
  OA22CHD U11726 ( .A1(n15369), .A2(n15416), .B1(n13339), .B2(n15236), .O(n15237) );
  OA22CHD U11727 ( .A1(n15106), .A2(n15416), .B1(n13339), .B2(n15120), .O(n15107) );
  OA22CHD U11728 ( .A1(n15015), .A2(n15416), .B1(n13339), .B2(n15014), .O(n15016) );
  OA22CHD U11729 ( .A1(n15043), .A2(n15416), .B1(n13339), .B2(n15042), .O(n15044) );
  ND2CHD U11730 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _87), .O(n14515) );
  OA22CHD U11731 ( .A1(n15040), .A2(n15420), .B1(n15047), .B2(n13339), .O(n14516) );
  ND2CHD U11732 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _94), .O(n14541) );
  OA22CHD U11733 ( .A1(n15035), .A2(n15420), .B1(n13339), .B2(n15046), .O(n14542) );
  ND2CHD U11734 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _101), .O(n14505) );
  OA22CHD U11735 ( .A1(n15352), .A2(n15420), .B1(n13339), .B2(n15040), .O(n14506) );
  ND2CHD U11736 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _108), .O(n14478) );
  OA22CHD U11737 ( .A1(n15029), .A2(n15420), .B1(n15035), .B2(n13339), .O(n14479) );
  ND2CHD U11738 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _115), .O(n14536) );
  OA22CHD U11739 ( .A1(n15337), .A2(n15416), .B1(n13339), .B2(n15348), .O(n15338) );
  OA22CHD U11740 ( .A1(n15488), .A2(n15416), .B1(n13339), .B2(n15349), .O(n15025) );
  OA22CHD U11741 ( .A1(n15345), .A2(n15416), .B1(n13339), .B2(n8982), .O(n15346) );
  OA22CHD U11742 ( .A1(n15030), .A2(n15416), .B1(n13339), .B2(n15050), .O(n15031) );
  OA22CHD U11743 ( .A1(n8982), .A2(n15420), .B1(n13339), .B2(n15036), .O(n15038) );
  ND2CHD U11744 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _44), .O(n14797) );
  ND2CHD U11745 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _51), .O(n14531) );
  OA22CHD U11746 ( .A1(n15036), .A2(n15420), .B1(n9528), .B2(n13339), .O(n14532) );
  OA22CHD U11747 ( .A1(n15286), .A2(n15416), .B1(n13339), .B2(n15285), .O(n15287) );
  ND2CHD U11748 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _97), .O(n15264) );
  OA22CHD U11749 ( .A1(n15386), .A2(n15416), .B1(n13339), .B2(n15284), .O(n13304) );
  ND2CHD U11750 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _61), .O(n14628) );
  OA22CHD U11751 ( .A1(n15293), .A2(n15420), .B1(n15064), .B2(n13339), .O(n14629) );
  ND2CHD U11752 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _125), .O(n15062) );
  ND2CHD U11753 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _86), .O(n15166) );
  ND2CHD U11754 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _93), .O(n14809) );
  ND2CHD U11755 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _100), .O(n15202) );
  ND2CHD U11756 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _107), .O(n15210) );
  ND2CHD U11757 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _114), .O(n15195) );
  OA22CHD U11758 ( .A1(n15461), .A2(n15416), .B1(n13339), .B2(n15214), .O(n13348) );
  OA22CHD U11759 ( .A1(n14904), .A2(n15416), .B1(n13339), .B2(n15198), .O(n14905) );
  ND2CHD U11760 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _57), .O(n15187) );
  ND2CHD U11761 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _121), .O(n14581) );
  OA22CHD U11762 ( .A1(n15189), .A2(n15420), .B1(n15209), .B2(n13339), .O(n14582) );
  OA22CHD U11763 ( .A1(n15462), .A2(n15416), .B1(n13339), .B2(n15205), .O(n14900) );
  OA22CHD U11764 ( .A1(n15130), .A2(n15416), .B1(n13339), .B2(n14817), .O(n13312) );
  OA22CHD U11765 ( .A1(n15317), .A2(n15416), .B1(n13339), .B2(n15169), .O(n13296) );
  OA22CHD U11766 ( .A1(n14814), .A2(n15416), .B1(n13339), .B2(n15172), .O(n14815) );
  OA22CHD U11767 ( .A1(n15169), .A2(n15420), .B1(n13339), .B2(n15185), .O(n14577) );
  ND2CHD U11768 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _36), .O(n14576) );
  OA22CHD U11769 ( .A1(n15120), .A2(n15420), .B1(n15089), .B2(n13339), .O(n14617) );
  ND2CHD U11770 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _48), .O(n14616) );
  ND2CHD U11771 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _55), .O(n14664) );
  OA22CHD U11772 ( .A1(n15128), .A2(n15420), .B1(n13339), .B2(n15092), .O(n14665) );
  ND2CHD U11773 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _62), .O(n15090) );
  ND2CHD U11774 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _117), .O(n14932) );
  ND2CHD U11775 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _110), .O(n14838) );
  ND2CHD U11776 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _103), .O(n14940) );
  ND2CHD U11777 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _96), .O(n14846) );
  OA22CHD U11778 ( .A1(n14924), .A2(n15416), .B1(n13339), .B2(n14923), .O(n14925) );
  OA22CHD U11779 ( .A1(n14919), .A2(n15420), .B1(n14931), .B2(n13339), .O(n14921) );
  ND2CHD U11780 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _60), .O(n14920) );
  ND2CHD U11781 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _124), .O(n14833) );
  OA22CHD U11782 ( .A1(n14321), .A2(n15416), .B1(n13339), .B2(n14943), .O(n13344) );
  OA22CHD U11783 ( .A1(n14302), .A2(n15416), .B1(n13339), .B2(n7392), .O(n13289) );
  OA22CHD U11784 ( .A1(n15452), .A2(n15416), .B1(n13339), .B2(n14957), .O(n14842) );
  OA22CHD U11785 ( .A1(n15483), .A2(n15416), .B1(n13339), .B2(n14945), .O(n14946) );
  OA22CHD U11786 ( .A1(n14802), .A2(n15416), .B1(n13339), .B2(n15150), .O(n13352) );
  OA22CHD U11787 ( .A1(n15055), .A2(n15416), .B1(n13339), .B2(n15413), .O(n15056) );
  OA22CHD U11788 ( .A1(n14866), .A2(n15416), .B1(n13339), .B2(n15423), .O(n14867) );
  OA22CHD U11789 ( .A1(n14880), .A2(n15416), .B1(n13339), .B2(n15421), .O(n14881) );
  OA22CHD U11790 ( .A1(n15141), .A2(n15416), .B1(n13339), .B2(n15140), .O(n15142) );
  OA22CHD U11791 ( .A1(n15426), .A2(n15420), .B1(n15146), .B2(n13339), .O(n15148) );
  OA22CHD U11792 ( .A1(n15393), .A2(n15416), .B1(n13339), .B2(n15404), .O(n15394) );
  OA22CHD U11793 ( .A1(n15400), .A2(n15416), .B1(n13339), .B2(n15399), .O(n15401) );
  ND2CHD U11794 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _49), .O(n14596) );
  OA22CHD U11795 ( .A1(n15404), .A2(n15420), .B1(n13339), .B2(n15296), .O(n14597) );
  ND2CHD U11796 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _56), .O(n15294) );
  ND2CHD U11797 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _63), .O(n14551) );
  OA22CHD U11798 ( .A1(n15296), .A2(n15420), .B1(n13339), .B2(n15426), .O(n14552) );
  ND2CHD U11799 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _127), .O(n15410) );
  OA22CHD U11800 ( .A1(n15417), .A2(n15416), .B1(n13339), .B2(n15415), .O(n15418) );
  OA22CHD U11801 ( .A1(n15075), .A2(n15416), .B1(n13339), .B2(n15074), .O(n15076) );
  ND2CHD U11802 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _88), .O(n14520) );
  ND2CHD U11803 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _102), .O(n14500) );
  ND2CHD U11804 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _123), .O(n15302) );
  ND2CHD U11805 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _59), .O(n15070) );
  OA22CHD U11806 ( .A1(n15069), .A2(n15420), .B1(n15304), .B2(n13339), .O(n15071) );
  ND2CHD U11807 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _45), .O(n14546) );
  OA22CHD U11808 ( .A1(n15224), .A2(n15416), .B1(n13339), .B2(n14557), .O(n13308) );
  XOR2EHD U11809 ( .I1(DOUT_18), .I2(n14103), .O(n13896) );
  ND2CHD U11810 ( .I1(n8189), .I2(n14412), .O(n14413) );
  OA12CHD U11811 ( .B1(n14709), .B2(n8189), .A1(n14708), .O(n14410) );
  ND2CHD U11812 ( .I1(n14713), .I2(n14414), .O(n14409) );
  ND2CHD U11813 ( .I1(n14688), .I2(n14680), .O(n14399) );
  OR2CHD U11814 ( .I1(n15243), .I2(n15422), .O(n14822) );
  OA112CHD U11815 ( .C1(n15420), .C2(n15247), .A1(n14821), .B1(n14820), .O(n14823) );
  ND2CHD U11816 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _91), .O(n14821) );
  OR2CHD U11817 ( .I1(n15340), .I2(n15422), .O(n13326) );
  OA112CHD U11818 ( .C1(n15420), .C2(n15014), .A1(n13325), .B1(n13324), .O(n13327) );
  ND2CHD U11819 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _2), .O(n13325) );
  NR2BHD U11820 ( .I1(n15254), .I2(n13277), .O(n14652) );
  NR2BHD U11821 ( .I1(n15285), .I2(n13277), .O(n14589) );
  OR2CHD U11822 ( .I1(n15289), .I2(n15422), .O(n14966) );
  OA112CHD U11823 ( .C1(n15420), .C2(n15281), .A1(n14965), .B1(n14964), .O(n14967) );
  ND2CHD U11824 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _76), .O(n14965) );
  OR2CHD U11825 ( .I1(n15280), .I2(n15422), .O(n15261) );
  OA112CHD U11826 ( .C1(n15420), .C2(n15277), .A1(n15260), .B1(n15259), .O(n15262) );
  ND2CHD U11827 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _90), .O(n15260) );
  OR2CHD U11828 ( .I1(n15267), .I2(n15422), .O(n14860) );
  ND2CHD U11829 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _26), .O(n14859) );
  OR2CHD U11830 ( .I1(n15191), .I2(n15422), .O(n15183) );
  OA112CHD U11831 ( .C1(n15420), .C2(n15182), .A1(n15181), .B1(n15180), .O(n15184) );
  ND2CHD U11832 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _72), .O(n15181) );
  AO12CHD U11833 ( .B1(n15367), .B2(n7043), .A1(n14899), .O(n6270) );
  ND2CHD U11834 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _50), .O(n14896) );
  OR2CHD U11835 ( .I1(n9478), .I2(n15422), .O(n14826) );
  OA112CHD U11836 ( .C1(n15420), .C2(n14954), .A1(n14825), .B1(n14824), .O(n14827) );
  ND2CHD U11837 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _82), .O(n14825) );
  OR2CHD U11838 ( .I1(n14927), .I2(n15422), .O(n14831) );
  ND2CHD U11839 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _68), .O(n14830) );
  ND2DHD U11840 ( .I1(n10174), .I2(n15139), .O(n6327) );
  NR2BHD U11841 ( .I1(n15421), .I2(n13277), .O(n14497) );
  OR2CHD U11842 ( .I1(n8662), .I2(n15422), .O(n14874) );
  ND2CHD U11843 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _28), .O(n14873) );
  OA112CHD U11844 ( .C1(n15422), .C2(n14991), .A1(n14990), .B1(n14989), .O(n14992) );
  OR2CHD U11845 ( .I1(n15306), .I2(n15422), .O(n13322) );
  OA112CHD U11846 ( .C1(n15420), .C2(n15073), .A1(n13321), .B1(n13320), .O(n13323) );
  ND2CHD U11847 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _67), .O(n13321) );
  OR2CHD U11848 ( .I1(n14976), .I2(n15422), .O(n14977) );
  ND2CHD U11849 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _81), .O(n14974) );
  NR2BHD U11850 ( .I1(n14483), .I2(n13277), .O(n14487) );
  OR2CHD U11851 ( .I1(n14499), .I2(n15422), .O(n13302) );
  OA112CHD U11852 ( .C1(n15420), .C2(n15074), .A1(n13301), .B1(n13300), .O(n13303) );
  ND2CHD U11853 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _17), .O(n13301) );
  ND2CHD U11854 ( .I1(n14465), .I2(_i_CLEFIA128_CON_T_x _2), .O(n14441) );
  NR2CHD U11855 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(_i_CLEFIA128_keyL _82), .O(n10561) );
  INVDHD U11856 ( .I(n10085), .O(n8576) );
  ND2DHD U11857 ( .I1(n9421), .I2(n7389), .O(n9420) );
  OA12EHD U11858 ( .B1(n8660), .B2(n8659), .A1(_i_CLEFIA128_state_reg _1), .O(n8658) );
  ND3CHD U11859 ( .I1(n8572), .I2(n8573), .I3(n7389), .O(n8571) );
  INVDHD U11860 ( .I(n11890), .O(n9932) );
  INVDHD U11861 ( .I(n10417), .O(n10199) );
  NR2CHD U11862 ( .I1(n9277), .I2(n9278), .O(n9908) );
  NR2EHD U11863 ( .I1(n15212), .I2(n9868), .O(n8735) );
  ND2DHD U11864 ( .I1(n8758), .I2(n12320), .O(n9813) );
  ND2DHD U11865 ( .I1(n12309), .I2(n12302), .O(n8540) );
  ND2HHD U11866 ( .I1(n8690), .I2(n6886), .O(n8689) );
  ND2CHD U11867 ( .I1(n9699), .I2(n12932), .O(n12933) );
  ND2DHD U11868 ( .I1(n12931), .I2(n10130), .O(n12932) );
  INVDHD U11869 ( .I(n12930), .O(n12931) );
  ND2HHD U11870 ( .I1(n12577), .I2(n12731), .O(n11089) );
  NR2BHD U11871 ( .I1(n11696), .I2(n8189), .O(n11698) );
  ND2CHD U11872 ( .I1(n6629), .I2(_i_CLEFIA128_keyK _118), .O(n11697) );
  ND3CHD U11873 ( .I1(n12596), .I2(n6990), .I3(n10376), .O(n10380) );
  ND2CHD U11874 ( .I1(n6846), .I2(n9648), .O(n10375) );
  ND2CHD U11875 ( .I1(n11648), .I2(n6837), .O(n11649) );
  ND2DHD U11876 ( .I1(n8962), .I2(n12869), .O(n10742) );
  ND2CHD U11877 ( .I1(n11440), .I2(n11192), .O(n10980) );
  ND2CHD U11878 ( .I1(n10978), .I2(n12450), .O(n10979) );
  ND2CHD U11879 ( .I1(n11178), .I2(n12501), .O(n10976) );
  ND3CHD U11880 ( .I1(n12479), .I2(n12464), .I3(n10974), .O(n10975) );
  NR2CHD U11881 ( .I1(n11939), .I2(n11938), .O(n9641) );
  ND2DHD U11882 ( .I1(n13459), .I2(n13439), .O(n11952) );
  ND2DHD U11883 ( .I1(n15353), .I2(_i_CLEFIA128_rndcnt_reg _0), .O(n11923) );
  NR2BHD U11884 ( .I1(n11914), .I2(n8189), .O(n11916) );
  ND2CHD U11885 ( .I1(n8224), .I2(_i_CLEFIA128_keyK _110), .O(n11915) );
  NR2CHD U11886 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(_i_CLEFIA128_keyK _110), .O(n11914) );
  INVGHD U11887 ( .I(n13024), .O(n12329) );
  ND2DHD U11888 ( .I1(n13442), .I2(n12422), .O(n10121) );
  ND2CHD U11889 ( .I1(n8185), .I2(n8223), .O(n13594) );
  NR2BHD U11890 ( .I1(n10573), .I2(n8189), .O(n10575) );
  ND2CHD U11891 ( .I1(n8224), .I2(_i_CLEFIA128_keyK _86), .O(n10574) );
  NR2CHD U11892 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(_i_CLEFIA128_keyK _86), .O(n10573) );
  ND2CHD U11893 ( .I1(n8215), .I2(n9348), .O(n12833) );
  ND2CHD U11894 ( .I1(n9559), .I2(n9348), .O(n10828) );
  INVCKGHD U11895 ( .I(n13084), .O(n11745) );
  ND2DHD U11896 ( .I1(n13550), .I2(n13513), .O(n12164) );
  ND2CHD U11897 ( .I1(n13366), .I2(n13028), .O(n13030) );
  ND2DHD U11898 ( .I1(n13570), .I2(_i_CLEFIA128_rndcnt_reg _0), .O(n11605) );
  NR2BHD U11899 ( .I1(n11602), .I2(n8189), .O(n11604) );
  ND2CHD U11900 ( .I1(n8224), .I2(_i_CLEFIA128_keyK _126), .O(n11603) );
  NR2CHD U11901 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(_i_CLEFIA128_keyK _126), .O(n11602) );
  ND2CHD U11902 ( .I1(n13194), .I2(n13187), .O(n12386) );
  ND2CHD U11903 ( .I1(n13024), .I2(n13373), .O(n12428) );
  ND2DHD U11904 ( .I1(n9283), .I2(n9693), .O(n9282) );
  MUX2CHD U11905 ( .A(n12017), .B(n12016), .S(_i_CLEFIA128_keyL _102), .O(n12022) );
  NR2BHD U11906 ( .I1(n12015), .I2(n8189), .O(n12017) );
  ND2CHD U11907 ( .I1(n6629), .I2(_i_CLEFIA128_keyK _102), .O(n12016) );
  NR2CHD U11908 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(_i_CLEFIA128_keyK _102), .O(n12015) );
  ND2CHD U11909 ( .I1(n8188), .I2(n7675), .O(n11359) );
  NR2CHD U11910 ( .I1(n9454), .I2(n10034), .O(n10811) );
  ND2CHD U11911 ( .I1(n12797), .I2(n12688), .O(n10812) );
  ND2DHD U11912 ( .I1(n13909), .I2(_i_CLEFIA128_rndcnt_reg _0), .O(n10338) );
  INVDHD U11913 ( .I(n8706), .O(n12929) );
  ND2CHD U11914 ( .I1(n11529), .I2(n11530), .O(n11449) );
  ND2CHD U11915 ( .I1(n11554), .I2(n6894), .O(n11445) );
  NR2BHD U11916 ( .I1(n11424), .I2(n11423), .O(n11425) );
  ND2CHD U11917 ( .I1(n13195), .I2(n13125), .O(n12006) );
  INVDHD U11918 ( .I(n14057), .O(n9578) );
  NR2CHD U11919 ( .I1(n13243), .I2(n9577), .O(n9576) );
  ND2DHD U11920 ( .I1(n8254), .I2(n8197), .O(n9577) );
  ND2CHD U11921 ( .I1(n13383), .I2(n13444), .O(n12222) );
  NR2CHD U11922 ( .I1(n9214), .I2(n12214), .O(n12215) );
  INVDHD U11923 ( .I(n13447), .O(n9233) );
  INVDHD U11924 ( .I(n12334), .O(n9588) );
  NR2BHD U11925 ( .I1(n12791), .I2(n12874), .O(n10970) );
  INVDHD U11926 ( .I(n8812), .O(n10950) );
  INVCKGHD U11927 ( .I(n10851), .O(n10136) );
  ND2DHD U11928 ( .I1(n12089), .I2(n11813), .O(n8842) );
  ND2CHD U11929 ( .I1(n8832), .I2(n11814), .O(n8843) );
  NR2CHD U11930 ( .I1(n13836), .I2(n12317), .O(n11791) );
  ND2CHD U11931 ( .I1(n12309), .I2(n12086), .O(n11733) );
  ND2CHD U11932 ( .I1(n11555), .I2(n11429), .O(n11431) );
  INVDHD U11933 ( .I(n12710), .O(n8963) );
  NR2CHD U11934 ( .I1(n7052), .I2(n12709), .O(n12711) );
  BUFJHD U11935 ( .I(n12681), .O(n9669) );
  ND2CHD U11936 ( .I1(n12376), .I2(n12268), .O(n12099) );
  ND3CHD U11937 ( .I1(n8393), .I2(n13122), .I3(n9886), .O(n9885) );
  ND2DHD U11938 ( .I1(n6589), .I2(n13099), .O(n13103) );
  NR2CHD U11939 ( .I1(n12808), .I2(n8912), .O(n12811) );
  MUX2CHD U11940 ( .A(n10489), .B(n10488), .S(_i_CLEFIA128_keyL _71), .O(n10494) );
  NR2BHD U11941 ( .I1(n10487), .I2(n8189), .O(n10489) );
  ND2CHD U11942 ( .I1(n8224), .I2(_i_CLEFIA128_keyK _71), .O(n10488) );
  NR2CHD U11943 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(_i_CLEFIA128_keyK _71), .O(n10487) );
  ND2CHD U11944 ( .I1(n11295), .I2(n11552), .O(n10997) );
  NR2EHD U11945 ( .I1(n10261), .I2(n12319), .O(n10260) );
  ND2CHD U11946 ( .I1(n13442), .I2(n8229), .O(n13443) );
  ND2DHD U11947 ( .I1(n13459), .I2(n13460), .O(n13462) );
  ND3CHD U11948 ( .I1(n13419), .I2(n13427), .I3(n13448), .O(n12243) );
  NR2CHD U11949 ( .I1(n13488), .I2(n13489), .O(n9365) );
  INVCKGHD U11950 ( .I(n13490), .O(n9375) );
  ND2HHD U11951 ( .I1(n11178), .I2(n12486), .O(n11432) );
  MUX2CHD U11952 ( .A(n10603), .B(n10602), .S(_i_CLEFIA128_keyL _87), .O(n10608) );
  NR2BHD U11953 ( .I1(n10601), .I2(n8189), .O(n10603) );
  ND2CHD U11954 ( .I1(n6629), .I2(_i_CLEFIA128_keyK _87), .O(n10602) );
  NR2CHD U11955 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(_i_CLEFIA128_keyK _87), .O(n10601) );
  NR2BHD U11956 ( .I1(n13388), .I2(n13422), .O(n13391) );
  ND3CHD U11957 ( .I1(n13024), .I2(n12350), .I3(n12426), .O(n11894) );
  ND2CHD U11958 ( .I1(n13134), .I2(n13629), .O(n13578) );
  ND2CHD U11959 ( .I1(n13573), .I2(n7031), .O(n13575) );
  ND3CHD U11960 ( .I1(n6918), .I2(n9463), .I3(n6897), .O(n13604) );
  NR2BHD U11961 ( .I1(n13619), .I2(n13618), .O(n13620) );
  ND2CHD U11962 ( .I1(n10713), .I2(n9047), .O(n10714) );
  NR2EHD U11963 ( .I1(n13461), .I2(n13017), .O(n9247) );
  ND2DHD U11964 ( .I1(n13603), .I2(n12280), .O(n9653) );
  ND2DHD U11965 ( .I1(n9006), .I2(n14055), .O(n12203) );
  NR2EHD U11966 ( .I1(n13210), .I2(n13209), .O(n13213) );
  ND2CHD U11967 ( .I1(n6529), .I2(n13589), .O(n13209) );
  ND3CHD U11968 ( .I1(n13596), .I2(n13194), .I3(n13164), .O(n12394) );
  ND2CHD U11969 ( .I1(n13183), .I2(n13182), .O(n13190) );
  NR2EHD U11970 ( .I1(n11488), .I2(n9417), .O(n9416) );
  NR2CHD U11971 ( .I1(n9467), .I2(n10894), .O(n10897) );
  ND2DHD U11972 ( .I1(n13790), .I2(_i_CLEFIA128_rndcnt_reg _0), .O(n10347) );
  ND2CHD U11973 ( .I1(n9625), .I2(n7705), .O(n11405) );
  NR2BHD U11974 ( .I1(n13578), .I2(n12921), .O(n12908) );
  NR2BHD U11975 ( .I1(n13152), .I2(n13176), .O(n12028) );
  ND2DHD U11976 ( .I1(n9003), .I2(n12674), .O(n10422) );
  ND2CHD U11977 ( .I1(n12743), .I2(n7705), .O(n11024) );
  ND3CHD U11978 ( .I1(n11042), .I2(n11371), .I3(n6956), .O(n11043) );
  NR2CHD U11979 ( .I1(n12977), .I2(n8681), .O(n12979) );
  NR2GHD U11980 ( .I1(n12102), .I2(n12101), .O(n12106) );
  NR2BHD U11981 ( .I1(n13645), .I2(n13644), .O(n13650) );
  ND2DHD U11982 ( .I1(n13651), .I2(n9210), .O(n13656) );
  ND3CHD U11983 ( .I1(n13653), .I2(n13652), .I3(n9309), .O(n13655) );
  ND2HHD U11984 ( .I1(n12324), .I2(n11959), .O(n13416) );
  ND3CHD U11985 ( .I1(n12283), .I2(n12285), .I3(n12284), .O(n12286) );
  NR2EHD U11986 ( .I1(n14139), .I2(n9161), .O(n9159) );
  ND2CHD U11987 ( .I1(n7017), .I2(KEY_3), .O(n13270) );
  NR2CHD U11988 ( .I1(n9173), .I2(n10924), .O(n8627) );
  INVDHD U11989 ( .I(n13278), .O(n10924) );
  ND2CHD U11990 ( .I1(n14682), .I2(n14681), .O(n14692) );
  ND2CHD U11991 ( .I1(n10928), .I2(DOUT_90), .O(n14699) );
  ND2CHD U11992 ( .I1(n10928), .I2(DOUT_24), .O(n13707) );
  ND2CHD U11993 ( .I1(n10928), .I2(DOUT_27), .O(n14149) );
  ND2CHD U11994 ( .I1(n10928), .I2(DOUT_28), .O(n14319) );
  ND2CHD U11995 ( .I1(n10928), .I2(DOUT_26), .O(n13875) );
  ND2CHD U11996 ( .I1(n10928), .I2(DOUT_15), .O(n14789) );
  ND2CHD U11997 ( .I1(n10928), .I2(DOUT_14), .O(n13956) );
  ND2CHD U11998 ( .I1(n10928), .I2(DOUT_13), .O(n15221) );
  ND2CHD U11999 ( .I1(n10928), .I2(DOUT_6), .O(n14021) );
  ND2CHD U12000 ( .I1(n10928), .I2(DOUT_4), .O(n10920) );
  ND2CHD U12001 ( .I1(n10928), .I2(DOUT_19), .O(n12820) );
  ND2CHD U12002 ( .I1(n10928), .I2(DOUT_93), .O(n14188) );
  ND2CHD U12003 ( .I1(n10928), .I2(DOUT_83), .O(n14371) );
  ND2CHD U12004 ( .I1(n10928), .I2(DOUT_5), .O(n14251) );
  OA22CHD U12005 ( .A1(n15400), .A2(n15513), .B1(n15512), .B2(n15055), .O(n13274) );
  ND2CHD U12006 ( .I1(n10928), .I2(DOUT_25), .O(n15459) );
  ND2CHD U12007 ( .I1(n10928), .I2(DOUT_10), .O(n13978) );
  ND2CHD U12008 ( .I1(n10928), .I2(DOUT_84), .O(n14381) );
  ND2CHD U12009 ( .I1(n10928), .I2(DOUT_81), .O(n14160) );
  ND2CHD U12010 ( .I1(n10928), .I2(DOUT_89), .O(n14889) );
  ND2CHD U12011 ( .I1(n10928), .I2(DOUT_91), .O(n14289) );
  ND2CHD U12012 ( .I1(n10928), .I2(DOUT_94), .O(n13694) );
  ND2CHD U12013 ( .I1(n10928), .I2(DOUT_95), .O(n14759) );
  ND2CHD U12014 ( .I1(n10928), .I2(DOUT_92), .O(n14279) );
  ND2CHD U12015 ( .I1(n10928), .I2(DOUT_85), .O(n14300) );
  ND2CHD U12016 ( .I1(n10928), .I2(DOUT_79), .O(n15358) );
  ND2CHD U12017 ( .I1(n10928), .I2(DOUT_87), .O(n13772) );
  ND2CHD U12018 ( .I1(n10928), .I2(DOUT_78), .O(n14035) );
  ND2CHD U12019 ( .I1(n10928), .I2(DOUT_8), .O(n15383) );
  ND2CHD U12020 ( .I1(n10928), .I2(DOUT_67), .O(n14336) );
  ND2CHD U12021 ( .I1(n10928), .I2(DOUT_88), .O(n14096) );
  ND2CHD U12022 ( .I1(n10928), .I2(DOUT_65), .O(n14235) );
  ND2CHD U12023 ( .I1(n10928), .I2(DOUT_86), .O(n13999) );
  ND2CHD U12024 ( .I1(n10928), .I2(DOUT_73), .O(n15005) );
  OA22CHD U12025 ( .A1(n15330), .A2(n15416), .B1(n13339), .B2(n15124), .O(n14820) );
  OA112CHD U12026 ( .C1(n15422), .C2(n15247), .A1(n15246), .B1(n15245), .O(n15248) );
  ND2CHD U12027 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _98), .O(n15245) );
  OA22CHD U12028 ( .A1(n15244), .A2(n15420), .B1(n15243), .B2(n13339), .O(n15246) );
  OA22CHD U12029 ( .A1(n15491), .A2(n15416), .B1(n13339), .B2(n15340), .O(n13316) );
  ND2CHD U12030 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _58), .O(n15020) );
  OR2CHD U12031 ( .I1(n9502), .I2(n13277), .O(n8449) );
  ND2CHD U12032 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _118), .O(n14586) );
  OA22CHD U12033 ( .A1(n15361), .A2(n15416), .B1(n13339), .B2(n15290), .O(n14964) );
  OA22CHD U12034 ( .A1(n15271), .A2(n15416), .B1(n13339), .B2(n15270), .O(n15272) );
  ND2CHD U12035 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _47), .O(n14961) );
  OA22CHD U12036 ( .A1(n15284), .A2(n15420), .B1(n13339), .B2(n15293), .O(n14962) );
  ND2CHD U12037 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _54), .O(n14659) );
  OA22CHD U12038 ( .A1(n15270), .A2(n15420), .B1(n13339), .B2(n15061), .O(n14660) );
  OA22CHD U12039 ( .A1(n15160), .A2(n15416), .B1(n13339), .B2(n15254), .O(n13336) );
  OA22CHD U12040 ( .A1(n15251), .A2(n15416), .B1(n13339), .B2(n15267), .O(n15252) );
  OA22CHD U12041 ( .A1(n14983), .A2(n15416), .B1(n13339), .B2(n15191), .O(n14984) );
  ND2CHD U12042 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _43), .O(n15173) );
  OA22CHD U12043 ( .A1(n15329), .A2(n15416), .B1(n13339), .B2(n15128), .O(n15111) );
  OA22CHD U12044 ( .A1(n15514), .A2(n15416), .B1(n13339), .B2(n14918), .O(n14850) );
  ND2CHD U12045 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _53), .O(n14622) );
  OA22CHD U12046 ( .A1(n14918), .A2(n15420), .B1(n13339), .B2(n14930), .O(n14623) );
  ND2CHD U12047 ( .I1(n10928), .I2(DOUT_75), .O(n14393) );
  ND2CHD U12048 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _85), .O(n14654) );
  OA22CHD U12049 ( .A1(n15137), .A2(n15420), .B1(n15058), .B2(n13339), .O(n14655) );
  ND2CHD U12050 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _99), .O(n14526) );
  OA22CHD U12051 ( .A1(n15146), .A2(n15420), .B1(n13339), .B2(n15407), .O(n14495) );
  ND2CHD U12052 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _113), .O(n14876) );
  OA22CHD U12053 ( .A1(n14608), .A2(n15416), .B1(n13339), .B2(n8662), .O(n13356) );
  ND2CHD U12054 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _116), .O(n14591) );
  ND2CHD U12055 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _95), .O(n14484) );
  OA22CHD U12056 ( .A1(n14291), .A2(n15416), .B1(n13339), .B2(n14499), .O(n13328) );
  ND2CHD U12057 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _52), .O(n14566) );
  OA22CHD U12058 ( .A1(n14972), .A2(n15420), .B1(n13339), .B2(n15301), .O(n14567) );
  OA22CHD U12059 ( .A1(n14979), .A2(n15420), .B1(n15069), .B2(n13339), .O(n14547) );
  ND2CHD U12060 ( .I1(n10928), .I2(DOUT_7), .O(n14777) );
  ND2CHD U12061 ( .I1(n10928), .I2(DOUT_72), .O(n14120) );
  OA22CHD U12062 ( .A1(n15428), .A2(n15416), .B1(n13339), .B2(n14979), .O(n13332) );
  NR2CHD U12063 ( .I1(n9173), .I2(n13278), .O(n13280) );
  NR2CHD U12064 ( .I1(n14444), .I2(n14678), .O(n13279) );
  ND2CHD U12065 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _38), .O(n14558) );
  OA22CHD U12066 ( .A1(n14557), .A2(n15420), .B1(n13339), .B2(n14972), .O(n14559) );
  ND2CHD U12067 ( .I1(n10928), .I2(DOUT_68), .O(n13259) );
  ND2CHD U12068 ( .I1(n10928), .I2(DOUT_0), .O(n15509) );
  OR2CHD U12069 ( .I1(_i_CLEFIA128_CON_T_xi _13), .I2(n14444), .O(n14445) );
  ND2CHD U12070 ( .I1(n14748), .I2(n7017), .O(n14725) );
  ND2CHD U12071 ( .I1(n14721), .I2(n14720), .O(n14722) );
  OR2CHD U12072 ( .I1(n15125), .I2(n15422), .O(n15126) );
  OA112CHD U12073 ( .C1(n15420), .C2(n15124), .A1(n15123), .B1(n15122), .O(n15127) );
  ND2CHD U12074 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _77), .O(n15123) );
  AO12CHD U12075 ( .B1(n15235), .B2(n7043), .A1(n15234), .O(n6335) );
  OA112CHD U12076 ( .C1(n15422), .C2(n15242), .A1(n15231), .B1(n15230), .O(n15232) );
  OA22CHD U12077 ( .A1(n9474), .A2(n15420), .B1(n15244), .B2(n13339), .O(n15231) );
  OR2CHD U12078 ( .I1(n15100), .I2(n15422), .O(n15087) );
  OA112CHD U12079 ( .C1(n15121), .C2(n15420), .A1(n15086), .B1(n15085), .O(n15088) );
  ND2CHD U12080 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _6), .O(n15086) );
  NR2BHD U12081 ( .I1(n15121), .I2(n13277), .O(n14513) );
  OR2CHD U12082 ( .I1(n15239), .I2(n15422), .O(n15104) );
  OA112CHD U12083 ( .C1(n15233), .C2(n15420), .A1(n15103), .B1(n15102), .O(n15105) );
  ND2CHD U12084 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _20), .O(n15103) );
  OR2CHD U12085 ( .I1(n15236), .I2(n15422), .O(n15109) );
  ND2CHD U12086 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _34), .O(n15108) );
  OR2CHD U12087 ( .I1(n15042), .I2(n15422), .O(n15018) );
  OA112CHD U12088 ( .C1(n15420), .C2(n15047), .A1(n15017), .B1(n15016), .O(n15019) );
  ND2CHD U12089 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _73), .O(n15017) );
  NR2BHD U12090 ( .I1(n8982), .I2(n13277), .O(n14518) );
  NR2BHD U12091 ( .I1(n15348), .I2(n13277), .O(n14508) );
  NR2BHD U12092 ( .I1(n15340), .I2(n13277), .O(n14539) );
  OR2CHD U12093 ( .I1(n15341), .I2(n15422), .O(n15342) );
  OA112CHD U12094 ( .C1(n15420), .C2(n15340), .A1(n15339), .B1(n15338), .O(n15343) );
  ND2CHD U12095 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _9), .O(n15339) );
  OR2CHD U12096 ( .I1(n15349), .I2(n15422), .O(n15350) );
  ND2CHD U12097 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _23), .O(n15347) );
  AO12CHD U12098 ( .B1(n7831), .B2(n7043), .A1(n15041), .O(n6255) );
  ND2CHD U12099 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _37), .O(n15037) );
  NR2BHD U12100 ( .I1(n15047), .I2(n13277), .O(n14534) );
  OR2CHD U12101 ( .I1(n15285), .I2(n15422), .O(n14856) );
  ND2CHD U12102 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _5), .O(n14855) );
  OR2CHD U12103 ( .I1(n15281), .I2(n15422), .O(n15282) );
  OA112CHD U12104 ( .C1(n15420), .C2(n15280), .A1(n15279), .B1(n15278), .O(n15283) );
  ND2CHD U12105 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _83), .O(n15279) );
  AO12CHD U12106 ( .B1(n15269), .B2(n7043), .A1(n15268), .O(n6322) );
  OA112CHD U12107 ( .C1(n15422), .C2(n15277), .A1(n15265), .B1(n15264), .O(n15266) );
  OA22CHD U12108 ( .A1(n15263), .A2(n15420), .B1(n15280), .B2(n13339), .O(n15265) );
  OR2CHD U12109 ( .I1(n15274), .I2(n15422), .O(n13306) );
  OA112CHD U12110 ( .C1(n15267), .C2(n15420), .A1(n13305), .B1(n13304), .O(n13307) );
  ND2CHD U12111 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _33), .O(n13305) );
  AO12CHD U12112 ( .B1(n15067), .B2(n7043), .A1(n15066), .O(n6280) );
  OA112CHD U12113 ( .C1(n15422), .C2(n15064), .A1(n15063), .B1(n15062), .O(n15065) );
  OA22CHD U12114 ( .A1(n15061), .A2(n15420), .B1(n15257), .B2(n13339), .O(n15063) );
  AO12CHD U12115 ( .B1(n15171), .B2(n7043), .A1(n15170), .O(n6320) );
  OA112CHD U12116 ( .C1(n15422), .C2(n15176), .A1(n15167), .B1(n15166), .O(n15168) );
  OA22CHD U12117 ( .A1(n15201), .A2(n15420), .B1(n15182), .B2(n13339), .O(n15167) );
  AO12CHD U12118 ( .B1(n15207), .B2(n7043), .A1(n15206), .O(n6333) );
  OA112CHD U12119 ( .C1(n15422), .C2(n15208), .A1(n15203), .B1(n15202), .O(n15204) );
  OA22CHD U12120 ( .A1(n15212), .A2(n15420), .B1(n13339), .B2(n15201), .O(n15203) );
  OA112CHD U12121 ( .C1(n15422), .C2(n15209), .A1(n15196), .B1(n15195), .O(n15197) );
  OA22CHD U12122 ( .A1(n15194), .A2(n15420), .B1(n15212), .B2(n13339), .O(n15196) );
  OR2CHD U12123 ( .I1(n15179), .I2(n15422), .O(n14907) );
  OA112CHD U12124 ( .C1(n15420), .C2(n15191), .A1(n14906), .B1(n14905), .O(n14908) );
  ND2CHD U12125 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _65), .O(n14906) );
  AO12CHD U12126 ( .B1(n15193), .B2(n7043), .A1(n15192), .O(n6277) );
  OA22CHD U12127 ( .A1(n15186), .A2(n15420), .B1(n13339), .B2(n15194), .O(n15188) );
  OR2CHD U12128 ( .I1(n15214), .I2(n15422), .O(n14902) );
  OA112CHD U12129 ( .C1(n15420), .C2(n15198), .A1(n14901), .B1(n14900), .O(n14903) );
  ND2CHD U12130 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _8), .O(n14901) );
  OR2CHD U12131 ( .I1(n14817), .I2(n15422), .O(n13298) );
  OA112CHD U12132 ( .C1(n15205), .C2(n15420), .A1(n13297), .B1(n13296), .O(n13299) );
  ND2CHD U12133 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _22), .O(n13297) );
  NR2BHD U12134 ( .I1(n15201), .I2(n13277), .O(n14579) );
  NR2BHD U12135 ( .I1(n15124), .I2(n13277), .O(n14667) );
  OA112CHD U12136 ( .C1(n15422), .C2(n14939), .A1(n14839), .B1(n14838), .O(n14840) );
  OA22CHD U12137 ( .A1(n14934), .A2(n15420), .B1(n14950), .B2(n13339), .O(n14839) );
  AO12CHD U12138 ( .B1(n15468), .B2(n7043), .A1(n14849), .O(n6323) );
  OA112CHD U12139 ( .C1(n15422), .C2(n14953), .A1(n14847), .B1(n14846), .O(n14848) );
  OA22CHD U12140 ( .A1(n15420), .A2(n14950), .B1(n14954), .B2(n13339), .O(n14847) );
  OR2CHD U12141 ( .I1(n7143), .I2(n15422), .O(n14916) );
  OA112CHD U12142 ( .C1(n9478), .C2(n15420), .A1(n14915), .B1(n14914), .O(n14917) );
  ND2CHD U12143 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _75), .O(n14915) );
  OR2CHD U12144 ( .I1(n14936), .I2(n15422), .O(n14928) );
  OA112CHD U12145 ( .C1(n15420), .C2(n14927), .A1(n14926), .B1(n14925), .O(n14929) );
  ND2CHD U12146 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _4), .O(n14926) );
  OA112CHD U12147 ( .C1(n15422), .C2(n14931), .A1(n14834), .B1(n14833), .O(n14835) );
  OA22CHD U12148 ( .A1(n14930), .A2(n15420), .B1(n14934), .B2(n13339), .O(n14834) );
  OR2CHD U12149 ( .I1(n14943), .I2(n15422), .O(n13294) );
  OA112CHD U12150 ( .C1(n14923), .C2(n15420), .A1(n13290), .B1(n13289), .O(n13295) );
  ND2CHD U12151 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _18), .O(n13290) );
  OR2CHD U12152 ( .I1(n14957), .I2(n15422), .O(n14948) );
  ND2CHD U12153 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _32), .O(n14947) );
  OR2CHD U12154 ( .I1(n15413), .I2(n15422), .O(n13354) );
  OA112CHD U12155 ( .C1(n15420), .C2(n15058), .A1(n13353), .B1(n13352), .O(n13355) );
  ND2CHD U12156 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _71), .O(n13353) );
  OR2CHD U12157 ( .I1(n15140), .I2(n15422), .O(n14883) );
  OA112CHD U12158 ( .C1(n15420), .C2(n15150), .A1(n14882), .B1(n14881), .O(n14884) );
  ND2CHD U12159 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _0), .O(n14882) );
  AO12CHD U12160 ( .B1(n15152), .B2(n7043), .A1(n15151), .O(n6285) );
  OA112CHD U12161 ( .C1(n15422), .C2(n15408), .A1(n15148), .B1(n15147), .O(n15149) );
  ND2CHD U12162 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _120), .O(n15147) );
  OR2CHD U12163 ( .I1(n15403), .I2(n15422), .O(n15396) );
  OA112CHD U12164 ( .C1(n15420), .C2(n8662), .A1(n15395), .B1(n15394), .O(n15397) );
  ND2CHD U12165 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _35), .O(n15395) );
  NR2BHD U12166 ( .I1(n15137), .I2(n13277), .O(n14599) );
  NR2BHD U12167 ( .I1(n15058), .I2(n13277), .O(n14554) );
  OR2CHD U12168 ( .I1(n15423), .I2(n15422), .O(n15424) );
  OA112CHD U12169 ( .C1(n15421), .C2(n15420), .A1(n15419), .B1(n15418), .O(n15425) );
  ND2CHD U12170 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _14), .O(n15419) );
  OR2CHD U12171 ( .I1(n15078), .I2(n15422), .O(n15079) );
  OA112CHD U12172 ( .C1(n15420), .C2(n15306), .A1(n15077), .B1(n15076), .O(n15080) );
  ND2CHD U12173 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _3), .O(n15077) );
  OR2CHD U12174 ( .I1(n15073), .I2(n15422), .O(n14970) );
  ND2CHD U12175 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _74), .O(n14969) );
  NR2BHD U12176 ( .I1(n14557), .I2(n13277), .O(n14523) );
  NR2BHD U12177 ( .I1(n14499), .I2(n13277), .O(n14503) );
  OA112CHD U12178 ( .C1(n15422), .C2(n15304), .A1(n15303), .B1(n15302), .O(n15305) );
  OA22CHD U12179 ( .A1(n15301), .A2(n15420), .B1(n15300), .B2(n13339), .O(n15303) );
  OR2CHD U12180 ( .I1(n14483), .I2(n15422), .O(n13310) );
  OA112CHD U12181 ( .C1(n15420), .C2(n14499), .A1(n13309), .B1(n13308), .O(n13311) );
  ND2CHD U12182 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _24), .O(n13309) );
  ND2CHD U12183 ( .I1(n14465), .I2(_i_CLEFIA128_CON_T_xi_2 ), .O(n14437) );
  MUXB2BHD U12184 ( .EB(n14744), .A(n14743), .B(n14742), .S(_i_CLEFIA128_CON_T_xi_2 ), .O(n14745) );
  MUX2CHD U12185 ( .A(n14738), .B(n14737), .S(_i_CLEFIA128_CON_T_x _6), .O(n14746) );
  NR2BHD U12186 ( .I1(n14733), .I2(n14748), .O(n14735) );
  NR2BHD U12187 ( .I1(n14732), .I2(n14432), .O(n14733) );
  NR2BHD U12188 ( .I1(n14728), .I2(n14748), .O(n14730) );
  ND2CHD U12189 ( .I1(n14465), .I2(_i_CLEFIA128_CON_T_xi _11), .O(n14461) );
  ND2CHD U12190 ( .I1(n14465), .I2(_i_CLEFIA128_CON_T_xi _13), .O(n14451) );
  NR2BHD U12191 ( .I1(n14412), .I2(n14709), .O(n14411) );
  NR2CHD U12192 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(_i_CLEFIA128_keyL _108), .O(n9272) );
  INVDHD U12193 ( .I(n11862), .O(n9273) );
  NR2GHD U12194 ( .I1(n10414), .I2(n14707), .O(n8930) );
  NR2CHD U12195 ( .I1(_i_CLEFIA128_keyL _44), .I2(n9989), .O(n9988) );
  ND2CHD U12196 ( .I1(n11575), .I2(n6851), .O(n11574) );
  INVDHD U12197 ( .I(n11668), .O(n8664) );
  NR2EHD U12198 ( .I1(n10544), .I2(n14707), .O(n10548) );
  ND2DHD U12199 ( .I1(n11891), .I2(n6851), .O(n10165) );
  ND2DHD U12200 ( .I1(n11891), .I2(n6851), .O(n10164) );
  ND2DHD U12201 ( .I1(n11675), .I2(n6851), .O(n10148) );
  ND2HHD U12202 ( .I1(n9132), .I2(_i_CLEFIA128_keyL _84), .O(n9131) );
  ND3CHD U12203 ( .I1(n10310), .I2(_i_CLEFIA128_rndcnt_reg _0), .I3(n15298), .O(n10311) );
  AN2HHD U12204 ( .I1(n8702), .I2(_i_CLEFIA128_state_reg _1), .O(n11988) );
  NR2EHD U12205 ( .I1(n9561), .I2(n10776), .O(n10025) );
  INVDHD U12206 ( .I(n7930), .O(n8697) );
  NR2BHD U12207 ( .I1(n13765), .I2(n7103), .O(n11690) );
  MUX2CHD U12208 ( .A(n11688), .B(n11687), .S(_i_CLEFIA128_keyL _119), .O(n11693) );
  NR2BHD U12209 ( .I1(n11686), .I2(n8189), .O(n11688) );
  ND2CHD U12210 ( .I1(n6629), .I2(_i_CLEFIA128_keyK _119), .O(n11687) );
  NR2CHD U12211 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(_i_CLEFIA128_keyK _119), .O(n11686) );
  ND2DHD U12212 ( .I1(n12309), .I2(n12299), .O(n8862) );
  ND2CHD U12213 ( .I1(n8224), .I2(_i_CLEFIA128_keyK _103), .O(n12008) );
  NR2BHD U12214 ( .I1(n12007), .I2(n8189), .O(n12009) );
  NR2CHD U12215 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(_i_CLEFIA128_keyK _103), .O(n12007) );
  NR2CHD U12216 ( .I1(n8969), .I2(n10444), .O(n8966) );
  ND2DHD U12217 ( .I1(n8564), .I2(n9916), .O(n10444) );
  INVGHD U12218 ( .I(n6842), .O(n10804) );
  NR2BHD U12219 ( .I1(n13995), .I2(n7103), .O(n11700) );
  ND2HHD U12220 ( .I1(n12192), .I2(n13084), .O(n11755) );
  INVGHD U12221 ( .I(n9367), .O(n13246) );
  MUX2CHD U12222 ( .A(n10499), .B(n10498), .S(_i_CLEFIA128_keyL _70), .O(n10502) );
  NR2BHD U12223 ( .I1(n10497), .I2(n8189), .O(n10499) );
  ND2CHD U12224 ( .I1(n8224), .I2(_i_CLEFIA128_keyK _70), .O(n10498) );
  NR2CHD U12225 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(_i_CLEFIA128_keyK _70), .O(n10497) );
  ND2DHD U12226 ( .I1(n9843), .I2(n11336), .O(n9842) );
  ND2DHD U12227 ( .I1(n13448), .I2(n9342), .O(n12245) );
  ND2CHD U12228 ( .I1(n13231), .I2(n7034), .O(n11848) );
  INVDHD U12229 ( .I(n13513), .O(n9153) );
  ND2CHD U12230 ( .I1(n8196), .I2(n10037), .O(n12065) );
  ND2DHD U12231 ( .I1(n13651), .I2(n9621), .O(n12090) );
  ND2CHD U12232 ( .I1(n10783), .I2(n10364), .O(n10365) );
  ND2DHD U12233 ( .I1(n14070), .I2(n13066), .O(n8648) );
  NR2CHD U12234 ( .I1(n8207), .I2(n6879), .O(n10435) );
  ND2CHD U12235 ( .I1(n11443), .I2(n11439), .O(n11001) );
  ND2DHD U12236 ( .I1(n11155), .I2(n11142), .O(n11144) );
  ND2CHD U12237 ( .I1(n12338), .I2(n13024), .O(n12339) );
  ND2DHD U12238 ( .I1(n12323), .I2(n13419), .O(n12326) );
  INVDHD U12239 ( .I(n8833), .O(n12351) );
  INVDHD U12240 ( .I(n9693), .O(n12966) );
  ND2CHD U12241 ( .I1(n11834), .I2(n11833), .O(n13234) );
  NR2BHD U12242 ( .I1(n11920), .I2(n8189), .O(n11922) );
  ND2CHD U12243 ( .I1(n8224), .I2(_i_CLEFIA128_keyK _111), .O(n11921) );
  NR2CHD U12244 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(_i_CLEFIA128_keyK _111), .O(n11920) );
  NR2BHD U12245 ( .I1(n14026), .I2(n6722), .O(n11918) );
  INVDHD U12246 ( .I(n12618), .O(n9259) );
  ND2HHD U12247 ( .I1(n9735), .I2(n10728), .O(n12875) );
  ND2DHD U12248 ( .I1(n9152), .I2(n13506), .O(n12146) );
  ND2HHD U12249 ( .I1(n9726), .I2(n12410), .O(n11931) );
  ND2CHD U12250 ( .I1(n13419), .I2(n13439), .O(n13034) );
  ND2CHD U12251 ( .I1(n10179), .I2(n12638), .O(n12639) );
  NR2BHD U12252 ( .I1(n13802), .I2(n7103), .O(n12019) );
  NR2CHD U12253 ( .I1(n13488), .I2(n11755), .O(n11632) );
  NR2EHD U12254 ( .I1(n8913), .I2(n8915), .O(n10823) );
  INVDHD U12255 ( .I(n8964), .O(n10822) );
  ND2CHD U12256 ( .I1(n13602), .I2(n13187), .O(n12047) );
  INVDHD U12257 ( .I(n9529), .O(n9514) );
  ND3CHD U12258 ( .I1(n6621), .I2(n10073), .I3(n8607), .O(n8609) );
  ND2DHD U12259 ( .I1(n8483), .I2(n11340), .O(n11110) );
  ND2CHD U12260 ( .I1(n8607), .I2(n11368), .O(n11109) );
  ND2CHD U12261 ( .I1(n13821), .I2(n13522), .O(n13523) );
  NR2EHD U12262 ( .I1(n12724), .I2(n10483), .O(n12556) );
  ND2CHD U12263 ( .I1(n9682), .I2(n12737), .O(n12583) );
  INVDHD U12264 ( .I(n9196), .O(n11463) );
  ND3CHD U12265 ( .I1(n8220), .I2(n11262), .I3(n11250), .O(n11084) );
  ND2CHD U12266 ( .I1(n12975), .I2(n7038), .O(n12976) );
  ND2DHD U12267 ( .I1(n13460), .I2(n13372), .O(n12984) );
  ND2DHD U12268 ( .I1(n13440), .I2(n12983), .O(n12985) );
  ND2DHD U12269 ( .I1(n12464), .I2(n12479), .O(n9140) );
  INVCHD U12270 ( .I(n11181), .O(n11182) );
  ND2CHD U12271 ( .I1(n11554), .I2(n11522), .O(n11149) );
  ND3CHD U12272 ( .I1(n12502), .I2(n12486), .I3(n9034), .O(n11148) );
  ND2HHD U12273 ( .I1(n12596), .I2(n10333), .O(n12648) );
  ND2DHD U12274 ( .I1(n6882), .I2(n10632), .O(n10333) );
  ND2CHD U12275 ( .I1(n6675), .I2(n12483), .O(n12485) );
  ND2CHD U12276 ( .I1(n8232), .I2(n7052), .O(n12701) );
  ND3CHD U12277 ( .I1(n14072), .I2(n13102), .I3(n14043), .O(n13089) );
  NR2BHD U12278 ( .I1(n11168), .I2(n11305), .O(n10571) );
  ND2CHD U12279 ( .I1(n12736), .I2(n12737), .O(n12739) );
  NR2CHD U12280 ( .I1(n14772), .I2(n7103), .O(n10491) );
  NR2BHD U12281 ( .I1(n10976), .I2(n10977), .O(n10982) );
  ND2CHD U12282 ( .I1(n11284), .I2(n12478), .O(n11008) );
  ND2CHD U12283 ( .I1(n11178), .I2(n12502), .O(n11004) );
  ND2CHD U12284 ( .I1(n12480), .I2(n11546), .O(n11550) );
  ND3CHD U12285 ( .I1(n12354), .I2(n12425), .I3(n13386), .O(n12355) );
  ND2DHD U12286 ( .I1(n13404), .I2(n11944), .O(n11945) );
  ND2CHD U12287 ( .I1(n13372), .I2(n12364), .O(n11947) );
  ND3CHD U12288 ( .I1(n13806), .I2(n8758), .I3(n13804), .O(n13807) );
  INVDHD U12289 ( .I(n13435), .O(n10094) );
  INVDHD U12290 ( .I(n13431), .O(n9213) );
  ND2DHD U12291 ( .I1(n13128), .I2(n12905), .O(n10221) );
  ND2CHD U12292 ( .I1(n11530), .I2(n10704), .O(n10705) );
  ND2CHD U12293 ( .I1(n11181), .I2(n9964), .O(n10696) );
  ND2CHD U12294 ( .I1(n9031), .I2(n10978), .O(n10688) );
  ND2CHD U12295 ( .I1(n11531), .I2(n12468), .O(n10689) );
  NR2CHD U12296 ( .I1(n13949), .I2(n7103), .O(n10393) );
  NR2BHD U12297 ( .I1(n10389), .I2(n8189), .O(n10391) );
  ND2CHD U12298 ( .I1(n8224), .I2(_i_CLEFIA128_keyK _78), .O(n10390) );
  NR2CHD U12299 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(_i_CLEFIA128_keyK _78), .O(n10389) );
  INVDHD U12300 ( .I(n8232), .O(n8513) );
  ND2CHD U12301 ( .I1(n6916), .I2(n12850), .O(n12852) );
  ND3CHD U12302 ( .I1(n9916), .I2(n7052), .I3(n12847), .O(n12848) );
  ND2DHD U12303 ( .I1(n6916), .I2(n12687), .O(n12700) );
  ND2CHD U12304 ( .I1(n10667), .I2(n12546), .O(n10686) );
  ND2CHD U12305 ( .I1(n10648), .I2(n9711), .O(n10655) );
  NR2EHD U12306 ( .I1(n9251), .I2(n13027), .O(n9250) );
  ND2CHD U12307 ( .I1(n14043), .I2(n14042), .O(n14045) );
  ND2DHD U12308 ( .I1(n12430), .I2(n13014), .O(n9286) );
  ND2CHD U12309 ( .I1(n12945), .I2(n12280), .O(n12282) );
  ND2CHD U12310 ( .I1(n13199), .I2(n13198), .O(n13202) );
  ND2CHD U12311 ( .I1(n6505), .I2(n13613), .O(n13197) );
  ND2CHD U12312 ( .I1(n9747), .I2(n13195), .O(n13196) );
  NR2CHD U12313 ( .I1(n9257), .I2(n11085), .O(n10878) );
  NR2CHD U12314 ( .I1(n12532), .I2(n12626), .O(n10840) );
  INVDHD U12315 ( .I(n7052), .O(n8507) );
  INVDHD U12316 ( .I(n10827), .O(n9854) );
  INVDHD U12317 ( .I(n8532), .O(n10814) );
  ND2DHD U12318 ( .I1(n9607), .I2(n7156), .O(n10475) );
  ND3CHD U12319 ( .I1(n12705), .I2(n12678), .I3(n8569), .O(n10887) );
  ND3CHD U12320 ( .I1(n8564), .I2(n8236), .I3(n8888), .O(n8570) );
  NR2BHD U12321 ( .I1(n13790), .I2(n6722), .O(n10348) );
  INVDHD U12322 ( .I(n6882), .O(n11222) );
  ND2DHD U12323 ( .I1(n9344), .I2(n12635), .O(n11223) );
  ND3CHD U12324 ( .I1(n9463), .I2(n12920), .I3(n13122), .O(n12922) );
  INVGHD U12325 ( .I(n7199), .O(n8751) );
  INVDHD U12326 ( .I(n12941), .O(n12942) );
  OR3EHD U12327 ( .I1(n11449), .I2(n11448), .I3(n11447), .O(n11450) );
  ND2CHD U12328 ( .I1(n11426), .I2(n11425), .O(n11427) );
  ND2DHD U12329 ( .I1(n8876), .I2(n12361), .O(n12244) );
  ND2DHD U12330 ( .I1(n13386), .I2(n9874), .O(n12249) );
  NR2CHD U12331 ( .I1(n9910), .I2(n12345), .O(n9909) );
  ND2CHD U12332 ( .I1(n12585), .I2(n11403), .O(n11121) );
  ND2CHD U12333 ( .I1(n11099), .I2(n11100), .O(n9534) );
  NR2CHD U12334 ( .I1(n10942), .I2(n8909), .O(n8953) );
  NR2CHD U12335 ( .I1(n11216), .I2(n11202), .O(n10287) );
  ND3CHD U12336 ( .I1(n12452), .I2(n12451), .I3(n12450), .O(n12461) );
  NR2BHD U12337 ( .I1(n12465), .I2(n12493), .O(n12466) );
  ND2DHD U12338 ( .I1(n12711), .I2(n9673), .O(n12712) );
  ND3CHD U12339 ( .I1(n12682), .I2(n9669), .I3(n8962), .O(n12684) );
  ND2CHD U12340 ( .I1(n9998), .I2(n12402), .O(n12112) );
  NR2CHD U12341 ( .I1(n9885), .I2(n12135), .O(n12136) );
  ND2DHD U12342 ( .I1(n8922), .I2(n12782), .O(n12786) );
  NR2EHD U12343 ( .I1(n9143), .I2(n8880), .O(n11524) );
  ND2DHD U12344 ( .I1(n13421), .I2(n13427), .O(n9337) );
  AN3EHD U12345 ( .I1(n13441), .I2(n13440), .I3(n13439), .O(n13453) );
  NR2CHD U12346 ( .I1(n9973), .I2(n13467), .O(n9113) );
  NR2CHD U12347 ( .I1(n10194), .I2(n9364), .O(n9363) );
  ND3CHD U12348 ( .I1(n11298), .I2(n9031), .I3(n11443), .O(n11299) );
  NR2CHD U12349 ( .I1(n13412), .I2(n13411), .O(n13414) );
  INVDHD U12350 ( .I(n13381), .O(n13395) );
  NR2CHD U12351 ( .I1(n13393), .I2(n13392), .O(n13394) );
  ND2CHD U12352 ( .I1(n13626), .I2(n13621), .O(n13586) );
  NR2BHD U12353 ( .I1(n13604), .I2(n13605), .O(n13606) );
  ND2CHD U12354 ( .I1(n13621), .I2(n13620), .O(n13623) );
  NR2BHD U12355 ( .I1(n8770), .I2(n11453), .O(n10717) );
  NR2BHD U12356 ( .I1(n10714), .I2(n11452), .O(n10715) );
  NR2BHD U12357 ( .I1(n12834), .I2(n12874), .O(n12835) );
  OR3EHD U12358 ( .I1(n12183), .I2(n12182), .I3(n13495), .O(n9069) );
  INVDHD U12359 ( .I(n13169), .O(n8715) );
  OR2EHD U12360 ( .I1(n13214), .I2(n10033), .O(n9769) );
  ND3CHD U12361 ( .I1(n11367), .I2(n11366), .I3(n9104), .O(n11373) );
  NR2BHD U12362 ( .I1(n8863), .I2(n11515), .O(n11408) );
  NR2BHD U12363 ( .I1(n12907), .I2(n12906), .O(n12909) );
  ND2CHD U12364 ( .I1(n10928), .I2(DOUT_21), .O(n14261) );
  ND2CHD U12365 ( .I1(n10928), .I2(DOUT_12), .O(n12890) );
  ND2CHD U12366 ( .I1(n10928), .I2(DOUT_66), .O(n15327) );
  ND2DHD U12367 ( .I1(n9173), .I2(BSY), .O(n13286) );
  ND2CHD U12368 ( .I1(n12996), .I2(n9947), .O(n12997) );
  BUFKHD U12369 ( .I(n14102), .O(n9761) );
  ND2CHD U12370 ( .I1(n10928), .I2(DOUT_31), .O(n13796) );
  ND2CHD U12371 ( .I1(n10928), .I2(DOUT_30), .O(n13917) );
  ND2CHD U12372 ( .I1(n10928), .I2(DOUT_29), .O(n15157) );
  ND2CHD U12373 ( .I1(n10928), .I2(DOUT_76), .O(n14310) );
  ND2CHD U12374 ( .I1(n10928), .I2(DOUT_23), .O(n13888) );
  ND2CHD U12375 ( .I1(n10928), .I2(DOUT_22), .O(n13990) );
  ND2CHD U12376 ( .I1(n10928), .I2(DOUT_17), .O(n13736) );
  ND2CHD U12377 ( .I1(n10928), .I2(DOUT_74), .O(n14356) );
  ND2CHD U12378 ( .I1(n10928), .I2(DOUT_18), .O(n13903) );
  ND2CHD U12379 ( .I1(n10928), .I2(DOUT_11), .O(n15314) );
  ND2CHD U12380 ( .I1(n10928), .I2(DOUT_1), .O(n13722) );
  OR2CHD U12381 ( .I1(n14384), .I2(n15512), .O(n10933) );
  AOI22BHD U12382 ( .A1(n7045), .A2(n9132), .B1(n15504), .B2(n10935), .O(n11128) );
  AO22CHD U12383 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _67), .B1(n15504), .B2(_i_CLEFIA128_keyK _3), .O(n13268) );
  ND2CHD U12384 ( .I1(n13292), .I2(n13269), .O(n13271) );
  ND2CHD U12385 ( .I1(n10928), .I2(DOUT_70), .O(n13856) );
  ND2CHD U12386 ( .I1(n10928), .I2(DOUT_69), .O(n14220) );
  AOI22BHD U12387 ( .A1(n7045), .A2(n15323), .B1(n15504), .B2(n15322), .O(n15335) );
  ND2CHD U12388 ( .I1(n10928), .I2(DOUT_16), .O(n13784) );
  ND2CHD U12389 ( .I1(n10928), .I2(DOUT_9), .O(n13759) );
  ND2CHD U12390 ( .I1(n10928), .I2(DOUT_82), .O(n13044) );
  ND2CHD U12391 ( .I1(n10928), .I2(DOUT_77), .O(n14206) );
  OA22CHD U12392 ( .A1(n14959), .A2(n15416), .B1(n13339), .B2(n15341), .O(n13324) );
  ND2CHD U12393 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _122), .O(n14637) );
  OA22CHD U12394 ( .A1(n14864), .A2(n15420), .B1(n15277), .B2(n13339), .O(n14650) );
  ND2CHD U12395 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _104), .O(n14649) );
  ND2CHD U12396 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _111), .O(n14862) );
  OA22CHD U12397 ( .A1(n15257), .A2(n15420), .B1(n15263), .B2(n13339), .O(n14863) );
  OA22CHD U12398 ( .A1(n15064), .A2(n15420), .B1(n14864), .B2(n13339), .O(n14587) );
  OA22CHD U12399 ( .A1(n15511), .A2(n15416), .B1(n13339), .B2(n9478), .O(n14951) );
  OA22CHD U12400 ( .A1(n15446), .A2(n15416), .B1(n13339), .B2(n14927), .O(n14914) );
  NR2BHD U12401 ( .I1(n8662), .I2(n13277), .O(n14657) );
  OA112CHD U12402 ( .C1(n15422), .C2(n15137), .A1(n15136), .B1(n15135), .O(n15138) );
  OA22CHD U12403 ( .A1(n15407), .A2(n15420), .B1(n15298), .B2(n13339), .O(n15136) );
  ND2CHD U12404 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _92), .O(n15135) );
  OA22CHD U12405 ( .A1(n15398), .A2(n15420), .B1(n15137), .B2(n13339), .O(n14527) );
  ND2CHD U12406 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _106), .O(n14494) );
  OA22CHD U12407 ( .A1(n14384), .A2(n15416), .B1(n13339), .B2(n15078), .O(n13320) );
  OA22CHD U12408 ( .A1(n14556), .A2(n15420), .B1(n13339), .B2(n14976), .O(n14521) );
  OA22CHD U12409 ( .A1(n14988), .A2(n15420), .B1(n13339), .B2(n14975), .O(n14485) );
  OA22CHD U12410 ( .A1(n14991), .A2(n15420), .B1(n14556), .B2(n13339), .O(n14501) );
  OA22CHD U12411 ( .A1(n14383), .A2(n15416), .B1(n13339), .B2(n14483), .O(n13300) );
  ND2CHD U12412 ( .I1(n10928), .I2(DOUT_71), .O(n15473) );
  ND2CHD U12413 ( .I1(n10928), .I2(DOUT_80), .O(n13943) );
  ND2CHD U12414 ( .I1(n10928), .I2(DOUT_2), .O(n13931) );
  ND2CHD U12415 ( .I1(n10928), .I2(DOUT_64), .O(n14130) );
  OA22CHD U12416 ( .A1(n14710), .A2(n14709), .B1(n8798), .B2(n14708), .O(n14712) );
  ND2CHD U12417 ( .I1(n14713), .I2(n14710), .O(n14711) );
  ND2CHD U12418 ( .I1(n14723), .I2(n15521), .O(n15523) );
  AOI22BHD U12419 ( .A1(n7045), .A2(n14362), .B1(n15504), .B2(n14361), .O(n14368) );
  ND2CHD U12420 ( .I1(n13983), .I2(n13982), .O(n6117) );
  AOI22BHD U12421 ( .A1(n7045), .A2(n14377), .B1(n15504), .B2(n14376), .O(n14378) );
  AOI22BHD U12422 ( .A1(n7045), .A2(n14275), .B1(n15504), .B2(n14274), .O(n14276) );
  ND2CHD U12423 ( .I1(n14240), .I2(n14239), .O(n6157) );
  AO12CHD U12424 ( .B1(n15440), .B2(n7043), .A1(n15101), .O(n6342) );
  OA112CHD U12425 ( .C1(n15422), .C2(n9474), .A1(n15098), .B1(n15097), .O(n15099) );
  OA22CHD U12426 ( .A1(n15096), .A2(n15420), .B1(n15242), .B2(n13339), .O(n15098) );
  OR2CHD U12427 ( .I1(n15121), .I2(n15422), .O(n13342) );
  OA112CHD U12428 ( .C1(n15420), .C2(n15125), .A1(n13341), .B1(n13340), .O(n13343) );
  ND2CHD U12429 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _70), .O(n13341) );
  OR2CHD U12430 ( .I1(n15233), .I2(n15422), .O(n15083) );
  ND2CHD U12431 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _13), .O(n15082) );
  OR2CHD U12432 ( .I1(n15249), .I2(n15422), .O(n15240) );
  ND2CHD U12433 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _27), .O(n15238) );
  OA12CHD U12434 ( .B1(n15499), .B2(n15106), .A1(n14997), .O(n14998) );
  OR2CHD U12435 ( .I1(n15047), .I2(n15422), .O(n15048) );
  ND2CHD U12436 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _80), .O(n15045) );
  NR2BHD U12437 ( .I1(n15349), .I2(n13277), .O(n14544) );
  NR2BHD U12438 ( .I1(n15341), .I2(n13277), .O(n14481) );
  OR2CHD U12439 ( .I1(n15014), .I2(n15422), .O(n13318) );
  ND2CHD U12440 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _66), .O(n13317) );
  OR2CHD U12441 ( .I1(n15348), .I2(n15422), .O(n15027) );
  ND2CHD U12442 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _16), .O(n15026) );
  OR2CHD U12443 ( .I1(n8982), .I2(n15422), .O(n15033) );
  OA112CHD U12444 ( .C1(n15420), .C2(n15349), .A1(n15032), .B1(n15031), .O(n15034) );
  ND2CHD U12445 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _30), .O(n15032) );
  AO12CHD U12446 ( .B1(n15435), .B2(n7043), .A1(n14800), .O(n6262) );
  OA22CHD U12447 ( .A1(n15050), .A2(n15420), .B1(n8902), .B2(n13339), .O(n14798) );
  AO12CHD U12448 ( .B1(n15024), .B2(n7043), .A1(n15023), .O(n6276) );
  OA112CHD U12449 ( .C1(n15422), .C2(n9528), .A1(n15021), .B1(n15020), .O(n15022) );
  OA22CHD U12450 ( .A1(n8902), .A2(n15420), .B1(n13339), .B2(n15344), .O(n15021) );
  OR2CHD U12451 ( .I1(n15284), .I2(n15422), .O(n15275) );
  ND2CHD U12452 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _40), .O(n15273) );
  NR2BHD U12453 ( .I1(n15281), .I2(n13277), .O(n14662) );
  NR2BHD U12454 ( .I1(n15289), .I2(n13277), .O(n14631) );
  OR2CHD U12455 ( .I1(n9502), .I2(n15422), .O(n8386) );
  OA112CHD U12456 ( .C1(n15420), .C2(n15285), .A1(n13337), .B1(n13336), .O(n13338) );
  ND2CHD U12457 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _12), .O(n13337) );
  OR2CHD U12458 ( .I1(n15254), .I2(n15422), .O(n15255) );
  ND2CHD U12459 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _19), .O(n15253) );
  OA12CHD U12460 ( .B1(n15499), .B2(n15251), .A1(n13361), .O(n13503) );
  OR2CHD U12461 ( .I1(n15182), .I2(n15422), .O(n14986) );
  OA112CHD U12462 ( .C1(n15420), .C2(n15176), .A1(n14985), .B1(n14984), .O(n14987) );
  ND2CHD U12463 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _79), .O(n14985) );
  AO12CHD U12464 ( .B1(n14813), .B2(n7043), .A1(n14812), .O(n6326) );
  OA22CHD U12465 ( .A1(n15208), .A2(n15420), .B1(n15176), .B2(n13339), .O(n14810) );
  AO12CHD U12466 ( .B1(n15392), .B2(n7043), .A1(n15215), .O(n6340) );
  OA112CHD U12467 ( .C1(n15422), .C2(n15212), .A1(n15211), .B1(n15210), .O(n15213) );
  OA22CHD U12468 ( .A1(n15209), .A2(n15420), .B1(n13339), .B2(n15208), .O(n15211) );
  OR2CHD U12469 ( .I1(n15198), .I2(n15422), .O(n13350) );
  OA112CHD U12470 ( .C1(n15420), .C2(n15179), .A1(n13349), .B1(n13348), .O(n13351) );
  ND2CHD U12471 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _1), .O(n13349) );
  NR2BHD U12472 ( .I1(n15179), .I2(n13277), .O(n14584) );
  OR2CHD U12473 ( .I1(n15205), .I2(n15422), .O(n13314) );
  ND2CHD U12474 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _15), .O(n13313) );
  OR2CHD U12475 ( .I1(n15169), .I2(n15422), .O(n14818) );
  OA112CHD U12476 ( .C1(n15420), .C2(n14817), .A1(n14816), .B1(n14815), .O(n14819) );
  ND2CHD U12477 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _29), .O(n14816) );
  AO12CHD U12478 ( .B1(n15178), .B2(n7043), .A1(n15177), .O(n6263) );
  OA22CHD U12479 ( .A1(n15172), .A2(n15420), .B1(n13339), .B2(n15186), .O(n15174) );
  OA12CHD U12480 ( .B1(n15499), .B2(n15271), .A1(n14980), .O(n14981) );
  ND2CHD U12481 ( .I1(n15200), .I2(n11130), .O(n14982) );
  OR2CHD U12482 ( .I1(n15120), .I2(n15422), .O(n15113) );
  ND2CHD U12483 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _41), .O(n15112) );
  NR2BHD U12484 ( .I1(n15243), .I2(n13277), .O(n14619) );
  OA22CHD U12485 ( .A1(n15089), .A2(n15420), .B1(n13339), .B2(n15096), .O(n15091) );
  OA12CHD U12486 ( .B1(n15499), .B2(n15130), .A1(n15129), .O(n15133) );
  AO12CHD U12487 ( .B1(n14938), .B2(n7043), .A1(n14937), .O(n6344) );
  OA112CHD U12488 ( .C1(n15422), .C2(n14934), .A1(n14933), .B1(n14932), .O(n14935) );
  OA22CHD U12489 ( .A1(n14931), .A2(n15420), .B1(n14939), .B2(n13339), .O(n14933) );
  AO12CHD U12490 ( .B1(n15131), .B2(n7043), .A1(n14944), .O(n6330) );
  OA112CHD U12491 ( .C1(n15422), .C2(n14950), .A1(n14941), .B1(n14940), .O(n14942) );
  OA22CHD U12492 ( .A1(n14939), .A2(n15420), .B1(n14953), .B2(n13339), .O(n14941) );
  OR2CHD U12493 ( .I1(n14923), .I2(n15422), .O(n13346) );
  OA112CHD U12494 ( .C1(n15420), .C2(n14936), .A1(n13345), .B1(n13344), .O(n13347) );
  ND2CHD U12495 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _11), .O(n13345) );
  OR2CHD U12496 ( .I1(n7392), .I2(n15422), .O(n14844) );
  ND2CHD U12497 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _25), .O(n14843) );
  OR2CHD U12498 ( .I1(n14945), .I2(n15422), .O(n14852) );
  OA112CHD U12499 ( .C1(n14957), .C2(n15420), .A1(n14851), .B1(n14850), .O(n14853) );
  ND2CHD U12500 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _39), .O(n14851) );
  AO12CHD U12501 ( .B1(n14913), .B2(n7043), .A1(n14912), .O(n6260) );
  ND2CHD U12502 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _46), .O(n14909) );
  NR2BHD U12503 ( .I1(n9478), .I2(n13277), .O(n14625) );
  OR2CHD U12504 ( .I1(n15058), .I2(n15422), .O(n15059) );
  OA112CHD U12505 ( .C1(n15420), .C2(n15298), .A1(n15057), .B1(n15056), .O(n15060) );
  ND2CHD U12506 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _78), .O(n15057) );
  OR2CHD U12507 ( .I1(n15421), .I2(n15422), .O(n14869) );
  OA112CHD U12508 ( .C1(n15420), .C2(n15140), .A1(n14868), .B1(n14867), .O(n14870) );
  ND2CHD U12509 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _7), .O(n14868) );
  OR2CHD U12510 ( .I1(n15150), .I2(n15422), .O(n15144) );
  OA112CHD U12511 ( .C1(n15413), .C2(n15420), .A1(n15143), .B1(n15142), .O(n15145) );
  ND2CHD U12512 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _64), .O(n15143) );
  AO12CHD U12513 ( .B1(n15520), .B2(n7043), .A1(n14879), .O(n6348) );
  OA112CHD U12514 ( .C1(n15422), .C2(n15146), .A1(n14877), .B1(n14876), .O(n14878) );
  OA22CHD U12515 ( .A1(n15408), .A2(n15420), .B1(n13339), .B2(n15398), .O(n14877) );
  OR2CHD U12516 ( .I1(n15404), .I2(n15422), .O(n15405) );
  ND2CHD U12517 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _42), .O(n15402) );
  AO12CHD U12518 ( .B1(n9817), .B2(n7043), .A1(n15299), .O(n6264) );
  OA22CHD U12519 ( .A1(n15399), .A2(n15420), .B1(n13339), .B2(n15409), .O(n15295) );
  AO12CHD U12520 ( .B1(n15481), .B2(n7043), .A1(n15414), .O(n6278) );
  OA22CHD U12521 ( .A1(n15409), .A2(n15420), .B1(n15408), .B2(n13339), .O(n15411) );
  OR2CHD U12522 ( .I1(n15415), .I2(n15422), .O(n13358) );
  ND2CHD U12523 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _21), .O(n13357) );
  NR2BHD U12524 ( .I1(n15078), .I2(n13277), .O(n14594) );
  OR2CHD U12525 ( .I1(n15074), .I2(n15422), .O(n13330) );
  OA112CHD U12526 ( .C1(n15420), .C2(n15078), .A1(n13329), .B1(n13328), .O(n13331) );
  ND2CHD U12527 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _10), .O(n13329) );
  NR2BHD U12528 ( .I1(n14976), .I2(n13277), .O(n14569) );
  NR2BHD U12529 ( .I1(n14975), .I2(n13277), .O(n14549) );
  OA12CHD U12530 ( .B1(n15499), .B2(n15475), .A1(n14769), .O(n14770) );
  OA12CHD U12531 ( .B1(n15499), .B2(n15400), .A1(n14672), .O(n14674) );
  ND2HHD U12532 ( .I1(n15193), .I2(n8257), .O(n9698) );
  OA12CHD U12533 ( .B1(n15499), .B2(n15115), .A1(n15012), .O(n15013) );
  OA12CHD U12534 ( .B1(n15499), .B2(n15369), .A1(n15368), .O(n15371) );
  OA12CHD U12535 ( .B1(n15499), .B2(n15373), .A1(n15372), .O(n15376) );
  OA12CHD U12536 ( .B1(n15499), .B2(n15437), .A1(n15436), .O(n15438) );
  ND2DHD U12537 ( .I1(n15367), .I2(n15500), .O(n8603) );
  OA12CHD U12538 ( .B1(n15499), .B2(n15360), .A1(n13962), .O(n13965) );
  OA12CHD U12539 ( .B1(n15499), .B2(n14302), .A1(n14172), .O(n14173) );
  OR2CHD U12540 ( .I1(n14557), .I2(n15422), .O(n13334) );
  ND2CHD U12541 ( .I1(n15504), .I2(_i_CLEFIA128_keyL _31), .O(n13333) );
  NR2BHD U12542 ( .I1(n14556), .I2(n13277), .O(n14561) );
  OA12CHD U12543 ( .B1(n15499), .B2(n15428), .A1(n15427), .O(n15429) );
  OA12CHD U12544 ( .B1(n15499), .B2(n15498), .A1(n15497), .O(n15502) );
  OA12CHD U12545 ( .B1(n15499), .B2(n15462), .A1(n13558), .O(n13559) );
  ND2CHD U12546 ( .I1(n15468), .I2(n11130), .O(n13561) );
  OA12CHD U12547 ( .B1(n14573), .B2(n15512), .A1(n14564), .O(n14565) );
  OA12CHD U12548 ( .B1(n8553), .B2(n15512), .A1(n8243), .O(n8217) );
  OA12CHD U12549 ( .B1(n15499), .B2(n15461), .A1(n13562), .O(n13563) );
  ND2CHD U12550 ( .I1(n15468), .I2(n15500), .O(n13565) );
  OA12CHD U12551 ( .B1(n15499), .B2(n15055), .A1(n14675), .O(n14677) );
  OA12CHD U12552 ( .B1(n15499), .B2(n15258), .A1(n15051), .O(n15052) );
  OA12CHD U12553 ( .B1(n15499), .B2(n14904), .A1(n14627), .O(n8244) );
  ND2DHD U12554 ( .I1(n15131), .I2(n15500), .O(n9729) );
  OA12CHD U12555 ( .B1(n15499), .B2(n15442), .A1(n15441), .O(n15443) );
  OA12CHD U12556 ( .B1(n15499), .B2(n15223), .A1(n14113), .O(n14114) );
  OA12CHD U12557 ( .B1(n15499), .B2(n14828), .A1(n14176), .O(n14177) );
  OA12CHD U12558 ( .B1(n15499), .B2(n15286), .A1(n13566), .O(n13568) );
  OA12CHD U12559 ( .B1(n15499), .B2(n15361), .A1(n13966), .O(n13968) );
  OA12CHD U12560 ( .B1(n15499), .B2(n15432), .A1(n15431), .O(n15433) );
  OA12CHD U12561 ( .B1(n15499), .B2(n15015), .A1(n14266), .O(n14267) );
  OA12CHD U12562 ( .B1(n15499), .B2(n15494), .A1(n15493), .O(n15496) );
  OA12EHD U12563 ( .B1(n14525), .B2(n15450), .A1(n8356), .O(n9856) );
  OA12CHD U12564 ( .B1(n15499), .B2(n15514), .A1(n13744), .O(n13745) );
  ND2CHD U12565 ( .I1(n15520), .I2(n11130), .O(n13747) );
  NR2BHD U12566 ( .I1(n14749), .I2(n14748), .O(n14751) );
  NR2BHD U12567 ( .I1(n14747), .I2(n14432), .O(n14749) );
  MUX2CHD U12568 ( .A(n14738), .B(n14737), .S(_i_CLEFIA128_CON_T_reg_4 ), .O(n14474) );
  ND2CHD U12569 ( .I1(n14465), .I2(_i_CLEFIA128_CON_T_x _7), .O(n14456) );
  ND2CHD U12570 ( .I1(n14465), .I2(_i_CLEFIA128_CON_T_x _10), .O(n14439) );
  MUX2CHD U12571 ( .A(n14738), .B(n14737), .S(_i_CLEFIA128_CON_T_x _12), .O(n14477) );
  MUX2CHD U12572 ( .A(n14738), .B(n14737), .S(_i_CLEFIA128_CON_T_x _14), .O(n14467) );
  MUX2CHD U12573 ( .A(n14738), .B(n14737), .S(_i_CLEFIA128_CON_T_x _0), .O(n14471) );
  MUX2CHD U12574 ( .A(n14708), .B(n14406), .S(n6851), .O(n14408) );
  MUX2CHD U12575 ( .A(n14423), .B(n14422), .S(_i_CLEFIA128_rndcnt_reg _4), .O(n14424) );
  ND2CHD U12576 ( .I1(n14418), .I2(_i_CLEFIA128_rndcnt_reg _3), .O(n14423) );
  AO12CHD U12577 ( .B1(n14713), .B2(n7048), .A1(_i_CLEFIA128_rndcnt_reg _2), .O(n14715) );
  ND2CHD U12578 ( .I1(n14726), .I2(_i_CLEFIA128_state_reg _0), .O(n14724) );
  MUX2CHD U12579 ( .A(_i_CLEFIA128_keyK _28), .B(KEY_28), .S(n7017), .O(n6375) );
  MUX2CHD U12580 ( .A(_i_CLEFIA128_keyK _27), .B(KEY_27), .S(n7017), .O(n6376) );
  MUX2CHD U12581 ( .A(_i_CLEFIA128_keyK _26), .B(KEY_26), .S(n7017), .O(n6377) );
  MUX2CHD U12582 ( .A(_i_CLEFIA128_keyK _25), .B(KEY_25), .S(n7017), .O(n6378) );
  MUX2CHD U12583 ( .A(_i_CLEFIA128_keyK _24), .B(KEY_24), .S(n7017), .O(n6379) );
  MUX2CHD U12584 ( .A(_i_CLEFIA128_keyK _23), .B(KEY_23), .S(n7017), .O(n6380) );
  MUX2CHD U12585 ( .A(_i_CLEFIA128_keyK _22), .B(KEY_22), .S(n7017), .O(n6381) );
  MUX2CHD U12586 ( .A(_i_CLEFIA128_keyK _21), .B(KEY_21), .S(n7017), .O(n6382) );
  MUX2CHD U12587 ( .A(_i_CLEFIA128_keyK _20), .B(KEY_20), .S(n7017), .O(n6383) );
  MUX2CHD U12588 ( .A(_i_CLEFIA128_keyK _19), .B(KEY_19), .S(n7017), .O(n6384) );
  MUX2CHD U12589 ( .A(_i_CLEFIA128_keyK _18), .B(KEY_18), .S(n7017), .O(n6385) );
  MUX2CHD U12590 ( .A(_i_CLEFIA128_keyK _17), .B(KEY_17), .S(n7017), .O(n6386) );
  MUX2CHD U12591 ( .A(_i_CLEFIA128_keyK _16), .B(KEY_16), .S(n7017), .O(n6387) );
  MUX2CHD U12592 ( .A(_i_CLEFIA128_keyK _15), .B(KEY_15), .S(n7017), .O(n6388) );
  MUX2CHD U12593 ( .A(_i_CLEFIA128_keyK _14), .B(KEY_14), .S(n7017), .O(n6389) );
  MUX2CHD U12594 ( .A(_i_CLEFIA128_keyK _13), .B(KEY_13), .S(n7017), .O(n6390) );
  MUX2CHD U12595 ( .A(_i_CLEFIA128_keyK _12), .B(KEY_12), .S(n7017), .O(n6391) );
  MUX2CHD U12596 ( .A(_i_CLEFIA128_keyK _11), .B(KEY_11), .S(n7017), .O(n6392) );
  MUX2CHD U12597 ( .A(_i_CLEFIA128_keyK _10), .B(KEY_10), .S(n7017), .O(n6393) );
  MUX2CHD U12598 ( .A(_i_CLEFIA128_keyK _9), .B(KEY_9), .S(n7017), .O(n6394));
  MUX2CHD U12599 ( .A(_i_CLEFIA128_keyK _8), .B(KEY_8), .S(n7017), .O(n6395));
  MUX2CHD U12600 ( .A(_i_CLEFIA128_keyK _7), .B(KEY_7), .S(n7017), .O(n6396));
  MUX2CHD U12601 ( .A(_i_CLEFIA128_keyK _6), .B(KEY_6), .S(n7017), .O(n6397));
  MUX2CHD U12602 ( .A(_i_CLEFIA128_keyK _5), .B(KEY_5), .S(n7017), .O(n6398));
  MUX2CHD U12603 ( .A(_i_CLEFIA128_keyK _4), .B(KEY_4), .S(n7017), .O(n6399));
  MUX2CHD U12604 ( .A(_i_CLEFIA128_keyK _3), .B(KEY_3), .S(n7017), .O(n6400));
  MUX2CHD U12605 ( .A(_i_CLEFIA128_keyK _2), .B(KEY_2), .S(n7017), .O(n6401));
  MUX2CHD U12606 ( .A(_i_CLEFIA128_keyK _1), .B(KEY_1), .S(n7017), .O(n6402));
  MUX2CHD U12607 ( .A(_i_CLEFIA128_keyK _127), .B(KEY_127), .S(n7017), .O(n6403) );
  MUX2CHD U12608 ( .A(_i_CLEFIA128_keyK _126), .B(KEY_126), .S(n7017), .O(n6404) );
  MUX2CHD U12609 ( .A(_i_CLEFIA128_keyK _125), .B(KEY_125), .S(n7017), .O(n6405) );
  MUX2CHD U12610 ( .A(_i_CLEFIA128_keyK _124), .B(KEY_124), .S(n7017), .O(n6406) );
  MUX2CHD U12611 ( .A(_i_CLEFIA128_keyK _123), .B(KEY_123), .S(n7017), .O(n6407) );
  MUX2CHD U12612 ( .A(_i_CLEFIA128_keyK _122), .B(KEY_122), .S(n7017), .O(n6408) );
  MUX2CHD U12613 ( .A(_i_CLEFIA128_keyK _121), .B(KEY_121), .S(n7017), .O(n6409) );
  MUX2CHD U12614 ( .A(_i_CLEFIA128_keyK _120), .B(KEY_120), .S(n7017), .O(n6410) );
  MUX2CHD U12615 ( .A(_i_CLEFIA128_keyK _119), .B(KEY_119), .S(n7017), .O(n6411) );
  MUX2CHD U12616 ( .A(_i_CLEFIA128_keyK _118), .B(KEY_118), .S(n7017), .O(n6412) );
  MUX2CHD U12617 ( .A(_i_CLEFIA128_keyK _117), .B(KEY_117), .S(n7017), .O(n6413) );
  MUX2CHD U12618 ( .A(_i_CLEFIA128_keyK _116), .B(KEY_116), .S(n7017), .O(n6414) );
  MUX2CHD U12619 ( .A(_i_CLEFIA128_keyK _115), .B(KEY_115), .S(n7017), .O(n6415) );
  MUX2CHD U12620 ( .A(_i_CLEFIA128_keyK _114), .B(KEY_114), .S(n7017), .O(n6416) );
  MUX2CHD U12621 ( .A(_i_CLEFIA128_keyK _113), .B(KEY_113), .S(n7017), .O(n6417) );
  MUX2CHD U12622 ( .A(_i_CLEFIA128_keyK _112), .B(KEY_112), .S(n7017), .O(n6418) );
  MUX2CHD U12623 ( .A(_i_CLEFIA128_keyK _111), .B(KEY_111), .S(n7017), .O(n6419) );
  MUX2CHD U12624 ( .A(_i_CLEFIA128_keyK _110), .B(KEY_110), .S(n7017), .O(n6420) );
  MUX2CHD U12625 ( .A(_i_CLEFIA128_keyK _109), .B(KEY_109), .S(n7017), .O(n6421) );
  MUX2CHD U12626 ( .A(_i_CLEFIA128_keyK _108), .B(KEY_108), .S(n7017), .O(n6422) );
  MUX2CHD U12627 ( .A(_i_CLEFIA128_keyK _107), .B(KEY_107), .S(n7017), .O(n6423) );
  MUX2CHD U12628 ( .A(_i_CLEFIA128_keyK _106), .B(KEY_106), .S(n7017), .O(n6424) );
  MUX2CHD U12629 ( .A(_i_CLEFIA128_keyK _105), .B(KEY_105), .S(n7017), .O(n6425) );
  MUX2CHD U12630 ( .A(_i_CLEFIA128_keyK _104), .B(KEY_104), .S(n7017), .O(n6426) );
  MUX2CHD U12631 ( .A(_i_CLEFIA128_keyK _103), .B(KEY_103), .S(n7017), .O(n6427) );
  MUX2CHD U12632 ( .A(_i_CLEFIA128_keyK _102), .B(KEY_102), .S(n7017), .O(n6428) );
  MUX2CHD U12633 ( .A(_i_CLEFIA128_keyK _101), .B(KEY_101), .S(n7017), .O(n6429) );
  MUX2CHD U12634 ( .A(_i_CLEFIA128_keyK _100), .B(KEY_100), .S(n7017), .O(n6430) );
  MUX2CHD U12635 ( .A(_i_CLEFIA128_keyK _99), .B(KEY_99), .S(n7017), .O(n6431) );
  MUX2CHD U12636 ( .A(_i_CLEFIA128_keyK _98), .B(KEY_98), .S(n7017), .O(n6432) );
  MUX2CHD U12637 ( .A(_i_CLEFIA128_keyK _97), .B(KEY_97), .S(n7017), .O(n6433) );
  MUX2CHD U12638 ( .A(_i_CLEFIA128_keyK _96), .B(KEY_96), .S(n7017), .O(n6434) );
  MUX2CHD U12639 ( .A(_i_CLEFIA128_keyK _95), .B(KEY_95), .S(n7017), .O(n6435) );
  MUX2CHD U12640 ( .A(_i_CLEFIA128_keyK _94), .B(KEY_94), .S(n7017), .O(n6436) );
  MUX2CHD U12641 ( .A(_i_CLEFIA128_keyK _93), .B(KEY_93), .S(n7017), .O(n6437) );
  MUX2CHD U12642 ( .A(_i_CLEFIA128_keyK _92), .B(KEY_92), .S(n7017), .O(n6438) );
  MUX2CHD U12643 ( .A(_i_CLEFIA128_keyK _91), .B(KEY_91), .S(n7017), .O(n6439) );
  MUX2CHD U12644 ( .A(_i_CLEFIA128_keyK _90), .B(KEY_90), .S(n7017), .O(n6440) );
  MUX2CHD U12645 ( .A(_i_CLEFIA128_keyK _89), .B(KEY_89), .S(n7017), .O(n6441) );
  MUX2CHD U12646 ( .A(_i_CLEFIA128_keyK _88), .B(KEY_88), .S(n7017), .O(n6442) );
  MUX2CHD U12647 ( .A(_i_CLEFIA128_keyK _87), .B(KEY_87), .S(n7017), .O(n6443) );
  MUX2CHD U12648 ( .A(_i_CLEFIA128_keyK _86), .B(KEY_86), .S(n7017), .O(n6444) );
  MUX2CHD U12649 ( .A(_i_CLEFIA128_keyK _85), .B(KEY_85), .S(n7017), .O(n6445) );
  MUX2CHD U12650 ( .A(_i_CLEFIA128_keyK _84), .B(KEY_84), .S(n7017), .O(n6446) );
  MUX2CHD U12651 ( .A(_i_CLEFIA128_keyK _83), .B(KEY_83), .S(n7017), .O(n6447) );
  MUX2CHD U12652 ( .A(_i_CLEFIA128_keyK _82), .B(KEY_82), .S(n7017), .O(n6448) );
  MUX2CHD U12653 ( .A(_i_CLEFIA128_keyK _81), .B(KEY_81), .S(n7017), .O(n6449) );
  MUX2CHD U12654 ( .A(_i_CLEFIA128_keyK _80), .B(KEY_80), .S(n7017), .O(n6450) );
  MUX2CHD U12655 ( .A(_i_CLEFIA128_keyK _79), .B(KEY_79), .S(n7017), .O(n6451) );
  MUX2CHD U12656 ( .A(_i_CLEFIA128_keyK _78), .B(KEY_78), .S(n7017), .O(n6452) );
  MUX2CHD U12657 ( .A(_i_CLEFIA128_keyK _77), .B(KEY_77), .S(n7017), .O(n6453) );
  MUX2CHD U12658 ( .A(_i_CLEFIA128_keyK _76), .B(KEY_76), .S(n7017), .O(n6454) );
  MUX2CHD U12659 ( .A(_i_CLEFIA128_keyK _75), .B(KEY_75), .S(n7017), .O(n6455) );
  MUX2CHD U12660 ( .A(_i_CLEFIA128_keyK _74), .B(KEY_74), .S(n7017), .O(n6456) );
  MUX2CHD U12661 ( .A(_i_CLEFIA128_keyK _73), .B(KEY_73), .S(n7017), .O(n6457) );
  MUX2CHD U12662 ( .A(_i_CLEFIA128_keyK _72), .B(KEY_72), .S(n7017), .O(n6458) );
  MUX2CHD U12663 ( .A(_i_CLEFIA128_keyK _71), .B(KEY_71), .S(n7017), .O(n6459) );
  MUX2CHD U12664 ( .A(_i_CLEFIA128_keyK _70), .B(KEY_70), .S(n7017), .O(n6460) );
  MUX2CHD U12665 ( .A(_i_CLEFIA128_keyK _69), .B(KEY_69), .S(n7017), .O(n6461) );
  MUX2CHD U12666 ( .A(_i_CLEFIA128_keyK _68), .B(KEY_68), .S(n7017), .O(n6462) );
  MUX2CHD U12667 ( .A(_i_CLEFIA128_keyK _67), .B(KEY_67), .S(n7017), .O(n6463) );
  MUX2CHD U12668 ( .A(_i_CLEFIA128_keyK _66), .B(KEY_66), .S(n7017), .O(n6464) );
  MUX2CHD U12669 ( .A(_i_CLEFIA128_keyK _65), .B(KEY_65), .S(n7017), .O(n6465) );
  MUX2CHD U12670 ( .A(_i_CLEFIA128_keyK _64), .B(KEY_64), .S(n7017), .O(n6466) );
  MUX2CHD U12671 ( .A(_i_CLEFIA128_keyK _63), .B(KEY_63), .S(n7017), .O(n6467) );
  MUX2CHD U12672 ( .A(_i_CLEFIA128_keyK _62), .B(KEY_62), .S(n7017), .O(n6468) );
  MUX2CHD U12673 ( .A(_i_CLEFIA128_keyK _61), .B(KEY_61), .S(n7017), .O(n6469) );
  MUX2CHD U12674 ( .A(_i_CLEFIA128_keyK _60), .B(KEY_60), .S(n7017), .O(n6470) );
  MUX2CHD U12675 ( .A(_i_CLEFIA128_keyK _59), .B(KEY_59), .S(n7017), .O(n6471) );
  MUX2CHD U12676 ( .A(_i_CLEFIA128_keyK _58), .B(KEY_58), .S(n7017), .O(n6472) );
  MUX2CHD U12677 ( .A(_i_CLEFIA128_keyK _57), .B(KEY_57), .S(n7017), .O(n6473) );
  MUX2CHD U12678 ( .A(_i_CLEFIA128_keyK _56), .B(KEY_56), .S(n7017), .O(n6474) );
  MUX2CHD U12679 ( .A(_i_CLEFIA128_keyK _55), .B(KEY_55), .S(n7017), .O(n6475) );
  MUX2CHD U12680 ( .A(_i_CLEFIA128_keyK _54), .B(KEY_54), .S(n7017), .O(n6476) );
  MUX2CHD U12681 ( .A(_i_CLEFIA128_keyK _53), .B(KEY_53), .S(n7017), .O(n6477) );
  MUX2CHD U12682 ( .A(_i_CLEFIA128_keyK _52), .B(KEY_52), .S(n7017), .O(n6478) );
  MUX2CHD U12683 ( .A(_i_CLEFIA128_keyK _51), .B(KEY_51), .S(n7017), .O(n6479) );
  MUX2CHD U12684 ( .A(_i_CLEFIA128_keyK _50), .B(KEY_50), .S(n7017), .O(n6480) );
  MUX2CHD U12685 ( .A(_i_CLEFIA128_keyK _49), .B(KEY_49), .S(n7017), .O(n6481) );
  MUX2CHD U12686 ( .A(_i_CLEFIA128_keyK _48), .B(KEY_48), .S(n7017), .O(n6482) );
  MUX2CHD U12687 ( .A(_i_CLEFIA128_keyK _47), .B(KEY_47), .S(n7017), .O(n6483) );
  MUX2CHD U12688 ( .A(_i_CLEFIA128_keyK _46), .B(KEY_46), .S(n7017), .O(n6484) );
  MUX2CHD U12689 ( .A(_i_CLEFIA128_keyK _45), .B(KEY_45), .S(n7017), .O(n6485) );
  MUX2CHD U12690 ( .A(_i_CLEFIA128_keyK _44), .B(KEY_44), .S(n7017), .O(n6486) );
  MUX2CHD U12691 ( .A(_i_CLEFIA128_keyK _43), .B(KEY_43), .S(n7017), .O(n6487) );
  MUX2CHD U12692 ( .A(_i_CLEFIA128_keyK _42), .B(KEY_42), .S(n7017), .O(n6488) );
  MUX2CHD U12693 ( .A(_i_CLEFIA128_keyK _41), .B(KEY_41), .S(n7017), .O(n6489) );
  MUX2CHD U12694 ( .A(_i_CLEFIA128_keyK _40), .B(KEY_40), .S(n7017), .O(n6490) );
  MUX2CHD U12695 ( .A(_i_CLEFIA128_keyK _39), .B(KEY_39), .S(n7017), .O(n6491) );
  MUX2CHD U12696 ( .A(_i_CLEFIA128_keyK _38), .B(KEY_38), .S(n7017), .O(n6492) );
  MUX2CHD U12697 ( .A(_i_CLEFIA128_keyK _37), .B(KEY_37), .S(n7017), .O(n6493) );
  MUX2CHD U12698 ( .A(_i_CLEFIA128_keyK _36), .B(KEY_36), .S(n7017), .O(n6494) );
  MUX2CHD U12699 ( .A(_i_CLEFIA128_keyK _35), .B(KEY_35), .S(n7017), .O(n6495) );
  MUX2CHD U12700 ( .A(_i_CLEFIA128_keyK _34), .B(KEY_34), .S(n7017), .O(n6496) );
  MUX2CHD U12701 ( .A(_i_CLEFIA128_keyK _33), .B(KEY_33), .S(n7017), .O(n6497) );
  MUX2CHD U12702 ( .A(_i_CLEFIA128_keyK _32), .B(KEY_32), .S(n7017), .O(n6498) );
  MUX2CHD U12703 ( .A(_i_CLEFIA128_keyK _31), .B(KEY_31), .S(n7017), .O(n6499) );
  MUX2CHD U12704 ( .A(_i_CLEFIA128_keyK _30), .B(KEY_30), .S(n7017), .O(n6500) );
  MUX2CHD U12705 ( .A(_i_CLEFIA128_keyK _29), .B(KEY_29), .S(n7017), .O(n6501) );
  MUX2CHD U12706 ( .A(_i_CLEFIA128_keyK _0), .B(KEY_0), .S(n7017), .O(n6502));
  AN2EHD U12707 ( .I1(n9129), .I2(n8801), .O(n8216) );
  AN2EHD U12708 ( .I1(n12975), .I2(n11904), .O(n8229) );
  INVGHD U12709 ( .I(n12989), .O(n9232) );
  AN3EHD U12710 ( .I1(n9529), .I2(n9631), .I3(n6571), .O(n8238) );
  INVDHD U12711 ( .I(n8606), .O(n9604) );
  AN2EHD U12712 ( .I1(n12448), .I2(n10615), .O(n8239) );
  AN3EHD U12713 ( .I1(n13684), .I2(n6582), .I3(n8736), .O(n8242) );
  AN2HHD U12714 ( .I1(n8454), .I2(n10534), .O(n8247) );
  AN2EHD U12715 ( .I1(n9230), .I2(n13487), .O(n8248) );
  NR3BHD U12716 ( .I1(n11442), .I2(n11441), .I3(n12493), .O(n8249) );
  INVDHD U12717 ( .I(n13478), .O(n11825) );
  AN2EHD U12718 ( .I1(n12487), .I2(n6894), .O(n8256) );
  INVDHD U12719 ( .I(n8547), .O(n10948) );
  AO22CHD U12720 ( .A1(n7045), .A2(n14116), .B1(n15504), .B2(n14115), .O(n8257) );
  AO22CHD U12721 ( .A1(n7045), .A2(n13950), .B1(n15504), .B2(n13949), .O(n8263) );
  AN2KHD U12722 ( .I1(n11959), .I2(n12335), .O(n8264) );
  OR2EHD U12723 ( .I1(n12082), .I2(n12318), .O(n8265) );
  AN3EHD U12724 ( .I1(n12928), .I2(n12040), .I3(n12041), .O(n8267) );
  AO22CHD U12725 ( .A1(n7045), .A2(n13571), .B1(n15504), .B2(n13570), .O(n8268) );
  AO22CHD U12726 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _110), .B1(n15504), .B2(_i_CLEFIA128_keyK _46), .O(n8269) );
  AO22CHD U12727 ( .A1(n7045), .A2(n13996), .B1(n15504), .B2(n13995), .O(n8270) );
  AO22CHD U12728 ( .A1(n7045), .A2(n13766), .B1(n15504), .B2(n13765), .O(n8271) );
  AO22CHD U12729 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _113), .B1(n15504), .B2(_i_CLEFIA128_keyK _49), .O(n8272) );
  AO22CHD U12730 ( .A1(n7045), .A2(n14202), .B1(n15504), .B2(n14201), .O(n8273) );
  AO22CHD U12731 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _125), .B1(n15504), .B2(_i_CLEFIA128_keyK _61), .O(n8274) );
  AO22CHD U12732 ( .A1(n7045), .A2(n14126), .B1(n15504), .B2(n14125), .O(n8275) );
  AO22CHD U12733 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _124), .B1(n15504), .B2(_i_CLEFIA128_keyK _60), .O(n8276) );
  AO22CHD U12734 ( .A1(n7045), .A2(n14012), .B1(n15504), .B2(n14011), .O(n8277) );
  AN2EHD U12735 ( .I1(n11485), .I2(n11510), .O(n8278) );
  AN2EHD U12736 ( .I1(n10051), .I2(n11679), .O(n8279) );
  AO22CHD U12737 ( .A1(n7045), .A2(n12827), .B1(n15504), .B2(n12826), .O(n8282) );
  AO22CHD U12738 ( .A1(n7045), .A2(n14326), .B1(n15504), .B2(n14325), .O(n8283) );
  AN3HHD U12739 ( .I1(n12192), .I2(n10296), .I3(n13479), .O(n8285) );
  AO22CHD U12740 ( .A1(n7045), .A2(n10304), .B1(n15504), .B2(n10303), .O(n8287) );
  AN2HHD U12741 ( .I1(n13018), .I2(n13420), .O(n8289) );
  AN2HHD U12742 ( .I1(n10122), .I2(n10121), .O(n8291) );
  AO22CHD U12743 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _84), .B1(n15504), .B2(_i_CLEFIA128_keyK _20), .O(n8293) );
  AO22CHD U12744 ( .A1(n7045), .A2(n14257), .B1(n15504), .B2(n14256), .O(n8295) );
  AN2EHD U12745 ( .I1(n11905), .I2(n9848), .O(n8296) );
  AO22CHD U12746 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _108), .B1(n15504), .B2(_i_CLEFIA128_keyK _44), .O(n8297) );
  INVDHD U12747 ( .I(n12840), .O(n9872) );
  OA12EHD U12748 ( .B1(n15499), .B2(n15317), .A1(n12142), .O(n8300) );
  AO22CHD U12749 ( .A1(n7045), .A2(n14307), .B1(n15504), .B2(n14306), .O(n8302) );
  AN2EHD U12750 ( .I1(n12323), .I2(n12439), .O(n8304) );
  AO22CHD U12751 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _92), .B1(n15504), .B2(_i_CLEFIA128_keyK _28), .O(n8306) );
  AN3EHD U12752 ( .I1(n11296), .I2(n11295), .I3(n9298), .O(n8308) );
  XNR2HHD U12753 ( .I1(_i_CLEFIA128_CON_T_x _3), .I2(DOUT_114), .O(n8310) );
  AO22CHD U12754 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _99), .B1(n15504), .B2(_i_CLEFIA128_keyK _35), .O(n8312) );
  OAI12CHD U12755 ( .B1(n15499), .B2(n15160), .A1(n14806), .O(n8313) );
  AN3EHD U12756 ( .I1(n13223), .I2(n7842), .I3(n10296), .O(n8316) );
  AN2EHD U12757 ( .I1(_i_CLEFIA128_keyK _10), .I2(_i_CLEFIA128_keyL _10), .O(n8317) );
  AN3EHD U12758 ( .I1(n11365), .I2(n11382), .I3(n11360), .O(n8318) );
  INVDHD U12759 ( .I(n9344), .O(n12528) );
  OR2KHD U12760 ( .I1(n9429), .I2(n12214), .O(n8320) );
  OR2HHD U12761 ( .I1(n12733), .I2(n12734), .O(n8321) );
  OR2EHD U12762 ( .I1(n12246), .I2(n12245), .O(n8322) );
  AN2EHD U12763 ( .I1(n8194), .I2(n8979), .O(n8323) );
  AN2EHD U12764 ( .I1(n13538), .I2(n9309), .O(n8325) );
  AN3EHD U12765 ( .I1(n13102), .I2(n8190), .I3(n13101), .O(n8326) );
  AN3EHD U12766 ( .I1(n13470), .I2(n9631), .I3(n13469), .O(n8327) );
  AN2EHD U12767 ( .I1(n11023), .I2(n12566), .O(n8330) );
  AN3HHD U12768 ( .I1(n9403), .I2(n14047), .I3(n14046), .O(n8332) );
  AN2EHD U12769 ( .I1(n12473), .I2(n12472), .O(n8335) );
  AN2EHD U12770 ( .I1(n6641), .I2(n8197), .O(n8336) );
  OR2EHD U12771 ( .I1(n9591), .I2(n9733), .O(n8339) );
  OR2KHD U12772 ( .I1(n8878), .I2(n9569), .O(n8340) );
  AN2HHD U12773 ( .I1(n8610), .I2(n13814), .O(n8341) );
  AN2HHD U12774 ( .I1(n10613), .I2(n10614), .O(n8343) );
  OR2EHD U12775 ( .I1(n10670), .I2(n7166), .O(n8344) );
  AN2EHD U12776 ( .I1(n11523), .I2(n10571), .O(n8347) );
  AN2EHD U12777 ( .I1(n13078), .I2(n13233), .O(n8348) );
  AN2EHD U12778 ( .I1(n13510), .I2(n13680), .O(n8351) );
  AN2EHD U12779 ( .I1(n12668), .I2(n10965), .O(n8352) );
  AN3HHD U12780 ( .I1(n9284), .I2(n8424), .I3(n12418), .O(n8353) );
  AN2EHD U12781 ( .I1(n9587), .I2(n9679), .O(n8357) );
  AN2EHD U12782 ( .I1(n10904), .I2(n10881), .O(n8359) );
  AN3HHD U12783 ( .I1(n14051), .I2(n13487), .I3(n14062), .O(n8362) );
  OAI13BHD U12784 ( .B1(n7199), .B2(n13206), .B3(n13205), .A1(n13608), .O(n8364) );
  INVDHD U12785 ( .I(_i_CLEFIA128_state_reg _1), .O(n8700) );
  AN3HHD U12786 ( .I1(n13824), .I2(n6684), .I3(n13819), .O(n8372) );
  AN2EHD U12787 ( .I1(n11875), .I2(_i_CLEFIA128_rndcnt_reg _0), .O(n8374) );
  AN3EHD U12788 ( .I1(n12013), .I2(n9477), .I3(_i_CLEFIA128_state_reg _1), .O(n8375) );
  AN3HHD U12789 ( .I1(n13596), .I2(n12402), .I3(n9603), .O(n8376) );
  AN2HHD U12790 ( .I1(n8812), .I2(n9003), .O(n8377) );
  XOR2EHD U12791 ( .I1(_i_CLEFIA128_CON_T_x _3), .I2(DOUT_50), .O(n8378) );
  AN2EHD U12792 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(_i_CLEFIA128_keyL _20), .O(n8381) );
  AN3HHD U12793 ( .I1(n11083), .I2(n11082), .I3(n12513), .O(n8382) );
  AN3EHD U12794 ( .I1(n8581), .I2(n9759), .I3(n13844), .O(n8384) );
  AOI22BHD U12795 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _78), .B1(n15504), .B2(_i_CLEFIA128_keyK _14), .O(n8388) );
  AOI22BHD U12796 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _118), .B1(n15504), .B2(_i_CLEFIA128_keyK _54), .O(n8389) );
  AN2HHD U12797 ( .I1(n9118), .I2(n9342), .O(n8392) );
  AN2EHD U12798 ( .I1(n12402), .I2(n9888), .O(n8393) );
  AN3EHD U12799 ( .I1(n13024), .I2(n13401), .I3(n9342), .O(n8394) );
  AN2EHD U12800 ( .I1(_i_CLEFIA128_keyK _29), .I2(_i_CLEFIA128_keyL _29), .O(n8396) );
  AN2HHD U12801 ( .I1(n12688), .I2(n12857), .O(n8398) );
  AN2EHD U12802 ( .I1(n12676), .I2(n8812), .O(n8399) );
  XOR2EHD U12803 ( .I1(_i_CLEFIA128_CON_T_xi _13), .I2(DOUT_126), .O(n8400));
  INVDHD U12804 ( .I(_i_CLEFIA128_state_reg _1), .O(n9989) );
  AN2EHD U12805 ( .I1(n12708), .I2(n12868), .O(n8403) );
  AN2EHD U12806 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(_i_CLEFIA128_keyL _16), .O(n8406) );
  AN2EHD U12807 ( .I1(n13439), .I2(n9574), .O(n8408) );
  AN2EHD U12808 ( .I1(n13600), .I2(n13601), .O(n8410) );
  AN2EHD U12809 ( .I1(n13550), .I2(n9210), .O(n8412) );
  INVDHD U12810 ( .I(n8495), .O(n12807) );
  AN3EHD U12811 ( .I1(n9916), .I2(n6670), .I3(n10207), .O(n8415) );
  AN2HHD U12812 ( .I1(n9355), .I2(n13482), .O(n8416) );
  AN3HHD U12813 ( .I1(n8472), .I2(n7025), .I3(n8318), .O(n8417) );
  ND2DHD U12814 ( .I1(n13592), .I2(n12945), .O(n8419) );
  AN3EHD U12815 ( .I1(n9806), .I2(n13085), .I3(n10296), .O(n8422) );
  AN2EHD U12816 ( .I1(n10966), .I2(n12858), .O(n8423) );
  ND2DHD U12817 ( .I1(n12422), .I2(n12423), .O(n8424) );
  ND2HHD U12818 ( .I1(n10421), .I2(n8921), .O(n12813) );
  AO22CHD U12819 ( .A1(n7045), .A2(n14316), .B1(n15504), .B2(n14315), .O(n8428) );
  AN2EHD U12820 ( .I1(n14864), .I2(_i_CLEFIA128_rndcnt_reg _0), .O(n8434) );
  AN2EHD U12821 ( .I1(n8901), .I2(n11661), .O(n8435) );
  AN2EHD U12822 ( .I1(_i_CLEFIA128_keyL _32), .I2(_i_CLEFIA128_keyK _32), .O(n8438) );
  OR2EHD U12823 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(_i_CLEFIA128_keyL _108), .O(n8439) );
  AN2HHD U12824 ( .I1(n10552), .I2(_i_CLEFIA128_state_reg _1), .O(n8440) );
  AN2EHD U12825 ( .I1(_i_CLEFIA128_keyK _18), .I2(_i_CLEFIA128_keyL _18), .O(n8445) );
  NR3BHD U12826 ( .I1(n12404), .I2(n13152), .I3(n12110), .O(n8446) );
  INVDHD U12827 ( .I(_i_CLEFIA128_keyL _6), .O(n9474) );
  OAI22CHD U12828 ( .A1(_i_CLEFIA128_keyK _3), .A2(n8222), .B1(n10300), .B2(_i_CLEFIA128_keyK _67), .O(n8450) );
  AN2HHD U12829 ( .I1(n8018), .I2(n11491), .O(n11371) );
  ND2CHD U12830 ( .I1(n8018), .I2(n11368), .O(n10509) );
  ND2HHD U12831 ( .I1(n8454), .I2(n12586), .O(n8453) );
  ND2CHD U12832 ( .I1(n8454), .I2(n12577), .O(n11035) );
  NR2GHD U12833 ( .I1(n8460), .I2(n8321), .O(n8459) );
  OAI12CHD U12834 ( .B1(n8468), .B2(n15416), .A1(n14595), .O(n6345) );
  OAI112BHD U12835 ( .C1(n8468), .C2(n15513), .A1(n14676), .B1(n14677), .O(n6161) );
  OAI112BHD U12836 ( .C1(n8468), .C2(n11129), .A1(n14673), .B1(n14674), .O(n6193) );
  ND3EHD U12837 ( .I1(n8465), .I2(n8467), .I3(n13276), .O(n6124) );
  XNR2KHD U12838 ( .I1(n9915), .I2(n9913), .O(n8468) );
  ND2HHD U12839 ( .I1(n8470), .I2(n12586), .O(n9353) );
  AN2CHD U12840 ( .I1(n8470), .I2(n11333), .O(n10513) );
  OA12HHD U12841 ( .B1(n8471), .B2(n11093), .A1(n12575), .O(n11108) );
  ND2HHD U12842 ( .I1(n8475), .I2(n8417), .O(n8471) );
  ND2HHD U12843 ( .I1(n8474), .I2(n9607), .O(n8473) );
  ND2KHD U12844 ( .I1(n12730), .I2(n11485), .O(n11409) );
  ND2HHD U12845 ( .I1(n8510), .I2(n11376), .O(n12759) );
  ND2HHD U12846 ( .I1(n9350), .I2(n12725), .O(n8477) );
  NR2CHD U12847 ( .I1(n12573), .I2(n11038), .O(n8478) );
  OR3HHD U12848 ( .I1(n8481), .I2(n11024), .I3(n11116), .O(n8480) );
  ND2HHD U12849 ( .I1(n10507), .I2(n8482), .O(n10508) );
  AN2HHD U12850 ( .I1(n7156), .I2(n12778), .O(n8482) );
  ND2HHD U12851 ( .I1(n9687), .I2(n7156), .O(n11397) );
  XOR2EHD U12852 ( .I1(n8486), .I2(DOUT_26), .O(n8550) );
  AN3HHD U12853 ( .I1(n8487), .I2(n11219), .I3(n11217), .O(n9573) );
  NR2GHD U12854 ( .I1(n10665), .I2(n9585), .O(n11219) );
  ND2HHD U12855 ( .I1(n9423), .I2(n12609), .O(n10665) );
  ND3EHD U12856 ( .I1(n8489), .I2(n8280), .I3(n8920), .O(n9382) );
  ND2HHD U12857 ( .I1(n8493), .I2(n8490), .O(n8725) );
  OR3HHD U12858 ( .I1(n10764), .I2(n9386), .I3(n8492), .O(n8491) );
  ND2CHD U12859 ( .I1(n8512), .I2(n8495), .O(n12843) );
  XOR2HHD U12860 ( .I1(_i_CLEFIA128_keyL _88), .I2(n8497), .O(n9421) );
  ND2HHD U12861 ( .I1(n6883), .I2(n9691), .O(n12598) );
  ND3EHD U12862 ( .I1(n8502), .I2(n10814), .I3(n8500), .O(n8499) );
  ND2HHD U12863 ( .I1(n10811), .I2(n12854), .O(n8501) );
  NR3BHD U12864 ( .I1(n10937), .I2(n8503), .I3(n8421), .O(n8502) );
  NR2GHD U12865 ( .I1(n10819), .I2(n8506), .O(n8505) );
  ND3EHD U12866 ( .I1(n12672), .I2(n10817), .I3(n10895), .O(n8506) );
  ND2KHD U12867 ( .I1(n9581), .I2(n10123), .O(n8508) );
  ND2HHD U12868 ( .I1(n8508), .I2(n8509), .O(n8532) );
  ND2KHD U12869 ( .I1(n7420), .I2(n7723), .O(n12677) );
  ND2KHD U12870 ( .I1(n9384), .I2(n8191), .O(n8511) );
  ND2CHD U12871 ( .I1(n12880), .I2(n8511), .O(n9386) );
  ND3EHD U12872 ( .I1(n8511), .I2(n8812), .I3(n12869), .O(n10439) );
  NR2BHD U12873 ( .I1(n12666), .I2(n8513), .O(n8512) );
  AN2CHD U12874 ( .I1(n8515), .I2(n11368), .O(n10533) );
  ND2HHD U12875 ( .I1(n8387), .I2(n8514), .O(n12721) );
  AN2EHD U12876 ( .I1(n8515), .I2(n7152), .O(n8514) );
  ND2KHD U12877 ( .I1(n8116), .I2(n7398), .O(n8515) );
  XOR2HHD U12878 ( .I1(n8516), .I2(n14246), .O(n10195) );
  XOR2HHD U12879 ( .I1(n9960), .I2(n8910), .O(n14246) );
  XOR2HHD U12880 ( .I1(n8517), .I2(n6798), .O(n8516) );
  XNR2KHD U12881 ( .I1(n9717), .I2(n9954), .O(n8519) );
  ND2HHD U12882 ( .I1(n8519), .I2(n8306), .O(n8518) );
  ND2KHD U12883 ( .I1(n8523), .I2(n8522), .O(n10259) );
  OAI12CHD U12884 ( .B1(n9008), .B2(n8530), .A1(n8529), .O(n8528) );
  ND3EHD U12885 ( .I1(n8546), .I2(n8545), .I3(n12690), .O(n9008) );
  NR2IHD U12886 ( .I1(n8533), .I2(n8694), .O(n8617) );
  ND2HHD U12887 ( .I1(n10466), .I2(n8369), .O(n10467) );
  NR2GHD U12888 ( .I1(n11396), .I2(n8534), .O(n11493) );
  ND3EHD U12889 ( .I1(n8535), .I2(n11482), .I3(n12729), .O(n8534) );
  AN2HHD U12890 ( .I1(n12089), .I2(n12088), .O(n13684) );
  INVCKGHD U12891 ( .I(n9067), .O(n12678) );
  NR2CHD U12892 ( .I1(n10947), .I2(n10944), .O(n8541) );
  NR2GHD U12893 ( .I1(n10937), .I2(n8542), .O(n12842) );
  OR2KHD U12894 ( .I1(n7886), .I2(n9067), .O(n10937) );
  NR2GHD U12895 ( .I1(n12808), .I2(n10936), .O(n10971) );
  XOR2HHD U12896 ( .I1(n8418), .I2(n13926), .O(n10196) );
  ND2KHD U12897 ( .I1(n9383), .I2(n8938), .O(n12690) );
  ND2KHD U12898 ( .I1(n10760), .I2(n9559), .O(n8888) );
  ND2KHD U12899 ( .I1(n9383), .I2(n8215), .O(n8962) );
  ND3EHD U12900 ( .I1(n8935), .I2(n8547), .I3(n12692), .O(n8934) );
  NR2GHD U12901 ( .I1(n10816), .I2(n10815), .O(n10895) );
  NR2IHD U12902 ( .I1(n9553), .I2(n9871), .O(n9378) );
  XNR3EHD U12903 ( .I1(n8793), .I2(n8550), .I3(n13895), .O(n8549) );
  OR2EHD U12904 ( .I1(n15513), .I2(n8553), .O(n10203) );
  OAI12CHD U12905 ( .B1(n8553), .B2(n15416), .A1(n8385), .O(n6338) );
  MUX2HHD U12906 ( .A(n13974), .B(n13975), .S(n8553), .O(n13983) );
  ND2KHD U12907 ( .I1(n10746), .I2(n9559), .O(n10888) );
  ND3EHD U12908 ( .I1(n8575), .I2(n8555), .I3(n8556), .O(n8554) );
  NR2EHD U12909 ( .I1(n10118), .I2(n8573), .O(n8555) );
  ND2HHD U12910 ( .I1(n8558), .I2(n8573), .O(n8557) );
  ND2HHD U12911 ( .I1(n8575), .I2(n8574), .O(n8558) );
  INVGHD U12912 ( .I(n8965), .O(n12687) );
  NR2IHD U12913 ( .I1(n10410), .I2(n14707), .O(n8560) );
  ND2HHD U12914 ( .I1(n9526), .I2(n8207), .O(n10428) );
  ND2KHD U12915 ( .I1(n12829), .I2(n8938), .O(n8564) );
  INVCKGHD U12916 ( .I(n8564), .O(n8593) );
  ND2HHD U12917 ( .I1(n8564), .I2(n10818), .O(n10820) );
  ND2HHD U12918 ( .I1(n10747), .I2(n8564), .O(n10957) );
  AN2HHD U12919 ( .I1(n8564), .I2(n8812), .O(n8565) );
  ND2HHD U12920 ( .I1(n14837), .I2(n11130), .O(n8566) );
  XNR2KHD U12921 ( .I1(_i_CLEFIA128_CON_T_xi_2 ), .I2(DOUT_43), .O(n8573) );
  ND2KHD U12922 ( .I1(n8899), .I2(n8346), .O(n8575) );
  ND2HHD U12923 ( .I1(n8579), .I2(n11774), .O(n11786) );
  ND2HHD U12924 ( .I1(n8581), .I2(n13805), .O(n8821) );
  ND3EHD U12925 ( .I1(n8581), .I2(n8655), .I3(n13510), .O(n8754) );
  ND2KHD U12926 ( .I1(n8209), .I2(n8178), .O(n8581) );
  AN2KHD U12927 ( .I1(n12312), .I2(n8583), .O(n13533) );
  XOR2HHD U12928 ( .I1(n14169), .I2(n14168), .O(n14805) );
  ND3EHD U12929 ( .I1(n9868), .I2(n15212), .I3(_i_CLEFIA128_rndcnt_reg _0), .O(n8587) );
  ND2KHD U12930 ( .I1(n8797), .I2(_i_CLEFIA128_keyK _8), .O(n9868) );
  ND2HHD U12931 ( .I1(n8590), .I2(_i_CLEFIA128_keyL _72), .O(n8588) );
  ND2HHD U12932 ( .I1(n8797), .I2(_i_CLEFIA128_keyK _72), .O(n8590) );
  ND2HHD U12933 ( .I1(n10964), .I2(n10966), .O(n8978) );
  INVNHD U12934 ( .I(n9857), .O(n9456) );
  ND2KHD U12935 ( .I1(n9320), .I2(n9317), .O(n9857) );
  OR3HHD U12936 ( .I1(n13172), .I2(n13574), .I3(n12097), .O(n8600) );
  ND3EHD U12937 ( .I1(n8891), .I2(n7009), .I3(n6529), .O(n8890) );
  XNR2KHD U12938 ( .I1(n13964), .I2(n8604), .O(n15367) );
  XOR2HHD U12939 ( .I1(n13963), .I2(n10139), .O(n8604) );
  ND3EHD U12940 ( .I1(n12905), .I2(n13602), .I3(n9127), .O(n12057) );
  NR2IHD U12941 ( .I1(n9037), .I2(n8606), .O(n8771) );
  ND2HHD U12942 ( .I1(n12719), .I2(n8608), .O(n11093) );
  ND2HHD U12943 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(_i_CLEFIA128_keyL _37), .O(n11973) );
  ND2HHD U12944 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(_i_CLEFIA128_keyL _53), .O(n9941) );
  ND2KHD U12945 ( .I1(n13132), .I2(n12915), .O(n8866) );
  ND2KHD U12946 ( .I1(n8196), .I2(n7036), .O(n13642) );
  NR2IHD U12947 ( .I1(n10026), .I2(n8611), .O(n13814) );
  ND3EHD U12948 ( .I1(n13493), .I2(n8613), .I3(n13228), .O(n10212) );
  ND2HHD U12949 ( .I1(n9433), .I2(n8614), .O(n9198) );
  ND2CHD U12950 ( .I1(n12835), .I2(n8615), .O(n12839) );
  OA13EHD U12951 ( .B1(n6533), .B2(n8620), .B3(n8619), .A1(n13826), .O(n8883));
  AN2HHD U12952 ( .I1(n8622), .I2(n10142), .O(n12091) );
  ND2KHD U12953 ( .I1(n12162), .I2(n13541), .O(n12300) );
  ND2HHD U12954 ( .I1(_i_CLEFIA128_keyL _52), .I2(_i_CLEFIA128_rndcnt_reg _0), .O(n9390) );
  OR3HHD U12955 ( .I1(n9236), .I2(n9068), .I3(n8624), .O(n9828) );
  OA13EHD U12956 ( .B1(n11738), .B2(n8624), .B3(n13657), .A1(n8294), .O(n9825));
  ND2KHD U12957 ( .I1(n12981), .I2(n12225), .O(n8625) );
  ND2KHD U12958 ( .I1(n10973), .I2(n10599), .O(n9208) );
  ND2HHD U12959 ( .I1(n9208), .I2(n8976), .O(n10120) );
  ND2HHD U12960 ( .I1(n9208), .I2(n9012), .O(n11447) );
  NR2GHD U12961 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(_i_CLEFIA128_keyL _117), .O(n8901) );
  INVCKGHD U12962 ( .I(_i_CLEFIA128_keyK _39), .O(n8626) );
  ND2HHD U12963 ( .I1(n8688), .I2(n8380), .O(n8687) );
  ND2HHD U12964 ( .I1(n10249), .I2(n8381), .O(n10248) );
  ND3EHD U12965 ( .I1(n10114), .I2(n15035), .I3(_i_CLEFIA128_rndcnt_reg _0), .O(n9205) );
  ND2CHD U12966 ( .I1(n6685), .I2(n8628), .O(n13648) );
  ND2KHD U12967 ( .I1(n8196), .I2(n7035), .O(n8628) );
  ND2HHD U12968 ( .I1(n8631), .I2(n8630), .O(n8629) );
  ND3EHD U12969 ( .I1(n9934), .I2(n10164), .I3(n11890), .O(n8630) );
  ND2HHD U12970 ( .I1(n9933), .I2(n9932), .O(n8631) );
  ND3EHD U12971 ( .I1(n9977), .I2(_i_CLEFIA128_rndcnt_reg _0), .I3(n14939), .O(n9976) );
  OA13EHD U12972 ( .B1(n11138), .B2(n8632), .B3(n11137), .A1(n12474), .O(n9045) );
  ND3EHD U12973 ( .I1(n10998), .I2(n10999), .I3(n11272), .O(n8632) );
  OAI12CHD U12974 ( .B1(n8980), .B2(n8639), .A1(n8563), .O(n8638) );
  ND3EHD U12975 ( .I1(n12672), .I2(n8640), .I3(n12792), .O(n8639) );
  ND3EHD U12976 ( .I1(n11581), .I2(n15078), .I3(_i_CLEFIA128_rndcnt_reg _0), .O(n11579) );
  ND2HHD U12977 ( .I1(n8644), .I2(n8642), .O(n9484) );
  NR2GHD U12978 ( .I1(n13494), .I2(n8646), .O(n8642) );
  ND2HHD U12979 ( .I1(n8326), .I2(n8647), .O(n8645) );
  XNR2KHD U12980 ( .I1(n9255), .I2(n9956), .O(n8651) );
  ND3CHD U12981 ( .I1(n6962), .I2(n12313), .I3(n8652), .O(n12096) );
  XOR2HHD U12982 ( .I1(_i_CLEFIA128_keyL _112), .I2(n11670), .O(n8653) );
  AN2CHD U12983 ( .I1(n8758), .I2(n8655), .O(n8654) );
  ND2KHD U12984 ( .I1(n7254), .I2(n7810), .O(n8655) );
  ND3EHD U12985 ( .I1(n13837), .I2(n13652), .I3(n8655), .O(n13507) );
  ND2CHD U12986 ( .I1(n8655), .I2(n13541), .O(n12155) );
  ND3EHD U12987 ( .I1(n8657), .I2(n10080), .I3(n13191), .O(n13605) );
  ND2CHD U12988 ( .I1(n9603), .I2(n8657), .O(n13146) );
  ND2HHD U12989 ( .I1(n8797), .I2(_i_CLEFIA128_keyK _49), .O(n11669) );
  ND2HHD U12990 ( .I1(n8661), .I2(n8658), .O(n8665) );
  ND3EHD U12991 ( .I1(n13474), .I2(n8327), .I3(n8666), .O(n13475) );
  NR3BHD U12992 ( .I1(n8668), .I2(n13473), .I3(n13472), .O(n8667) );
  ND2HHD U12993 ( .I1(n8669), .I2(n8264), .O(n10182) );
  ND3EHD U12994 ( .I1(n8674), .I2(n8671), .I3(n8670), .O(n8669) );
  NR3BHD U12995 ( .I1(n12244), .I2(n9439), .I3(n13376), .O(n8674) );
  ND3EHD U12996 ( .I1(n8429), .I2(n8677), .I3(n8676), .O(n8675) );
  OR3HHD U12997 ( .I1(n9973), .I2(n8681), .I3(n11958), .O(n11960) );
  OR3HHD U12998 ( .I1(n11954), .I2(n11955), .I3(n12440), .O(n8681) );
  ND2HHD U12999 ( .I1(n12554), .I2(n12555), .O(n12746) );
  ND2HHD U13000 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(_i_CLEFIA128_keyL _59), .O(n11580) );
  ND2HHD U13001 ( .I1(n10545), .I2(n8370), .O(n10546) );
  ND3CHD U13002 ( .I1(n8685), .I2(n12863), .I3(n12862), .O(n12865) );
  ND2KHD U13003 ( .I1(n8908), .I2(n9383), .O(n12880) );
  NR2CHD U13004 ( .I1(n8963), .I2(n8686), .O(n9673) );
  NR2EHD U13005 ( .I1(n8686), .I2(n8809), .O(n8807) );
  ND2HHD U13006 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(_i_CLEFIA128_keyL _41), .O(n11880) );
  ND3EHD U13007 ( .I1(n10553), .I2(n15244), .I3(_i_CLEFIA128_rndcnt_reg _0), .O(n10552) );
  ND3EHD U13008 ( .I1(n10456), .I2(_i_CLEFIA128_rndcnt_reg _0), .I3(n14934), .O(n10457) );
  ND3EHD U13009 ( .I1(n10461), .I2(_i_CLEFIA128_rndcnt_reg _0), .I3(n15209), .O(n10462) );
  ND3EHD U13010 ( .I1(n11672), .I2(_i_CLEFIA128_rndcnt_reg _0), .I3(n15179), .O(n11673) );
  ND2HHD U13011 ( .I1(n12163), .I2(n9808), .O(n8693) );
  ND3EHD U13012 ( .I1(n13652), .I2(n8695), .I3(n13671), .O(n8694) );
  ND2HHD U13013 ( .I1(n8696), .I2(n8178), .O(n8695) );
  NR2GHD U13014 ( .I1(n8700), .I2(n8699), .O(n8698) );
  OAI12CHD U13015 ( .B1(n8705), .B2(n15416), .A1(n8360), .O(n6282) );
  NR2IHD U13016 ( .I1(n8713), .I2(n8707), .O(n14106) );
  ND3EHD U13017 ( .I1(n8709), .I2(n8708), .I3(n8364), .O(n8707) );
  OAI12CHD U13018 ( .B1(n9878), .B2(n9769), .A1(n13585), .O(n8708) );
  XOR2HHD U13019 ( .I1(n9592), .I2(n14106), .O(n14107) );
  ND3EHD U13020 ( .I1(n8712), .I2(n8711), .I3(n13180), .O(n8710) );
  OA12HHD U13021 ( .B1(n9629), .B2(n8714), .A1(n13634), .O(n8713) );
  XOR2HHD U13022 ( .I1(n13779), .I2(n9893), .O(n15374) );
  NR2GHD U13023 ( .I1(n9728), .I2(n8716), .O(n9727) );
  ND3EHD U13024 ( .I1(n7011), .I2(n12928), .I3(n10186), .O(n8716) );
  OAI12CHD U13025 ( .B1(n12383), .B2(n12902), .A1(n11995), .O(n12124) );
  NR2GHD U13026 ( .I1(n7023), .I2(n8815), .O(n12304) );
  XOR2HHD U13027 ( .I1(n13701), .I2(n8719), .O(n14143) );
  XOR2HHD U13028 ( .I1(n14102), .I2(n10017), .O(n10229) );
  ND3EHD U13029 ( .I1(n11078), .I2(n10790), .I3(n12545), .O(n8720) );
  ND3EHD U13030 ( .I1(n10780), .I2(n12516), .I3(n12650), .O(n8721) );
  ND3EHD U13031 ( .I1(n8726), .I2(n8724), .I3(n8722), .O(n14102) );
  ND2HHD U13032 ( .I1(n8725), .I2(n12671), .O(n8724) );
  ND3EHD U13033 ( .I1(n8727), .I2(n8728), .I3(n12717), .O(n8726) );
  ND3EHD U13034 ( .I1(n9381), .I2(n9380), .I3(n8231), .O(n8727) );
  ND3EHD U13035 ( .I1(n9638), .I2(n9379), .I3(n12805), .O(n8728) );
  ND3EHD U13036 ( .I1(n9127), .I2(n12390), .I3(n8729), .O(n13114) );
  ND2CHD U13037 ( .I1(n9012), .I2(n12450), .O(n11007) );
  ND2KHD U13038 ( .I1(n9800), .I2(n7671), .O(n9012) );
  ND2KHD U13039 ( .I1(n9359), .I2(n10588), .O(n11452) );
  ND2HHD U13040 ( .I1(n12453), .I2(n6764), .O(n11139) );
  ND2KHD U13041 ( .I1(n9800), .I2(n10600), .O(n9359) );
  ND3EHD U13042 ( .I1(n8731), .I2(n8733), .I3(n14314), .O(n6146) );
  ND2HHD U13043 ( .I1(n8732), .I2(n8297), .O(n8731) );
  INVGHD U13044 ( .I(n8734), .O(n8732) );
  XOR2HHD U13045 ( .I1(n10019), .I2(n10020), .O(n8734) );
  OA13EHD U13046 ( .B1(n12391), .B2(n12392), .B3(n8737), .A1(n13622), .O(n9860) );
  NR2GHD U13047 ( .I1(n10157), .I2(n15191), .O(n8738) );
  ND2CHD U13048 ( .I1(n9084), .I2(n13398), .O(n11900) );
  ND2KHD U13049 ( .I1(n12423), .I2(n7032), .O(n9084) );
  ND2HHD U13050 ( .I1(n11986), .I2(n8740), .O(n9321) );
  NR2GHD U13051 ( .I1(n15257), .I2(n9789), .O(n8743) );
  AN2HHD U13052 ( .I1(n12029), .I2(n12001), .O(n9189) );
  XNR2KHD U13053 ( .I1(n11969), .I2(n8747), .O(n12029) );
  XOR2HHD U13054 ( .I1(n8749), .I2(n8748), .O(n14813) );
  XOR2HHD U13055 ( .I1(n13360), .I2(n14014), .O(n8748) );
  XOR2HHD U13056 ( .I1(n14016), .I2(n13912), .O(n8749) );
  ND3EHD U13057 ( .I1(n7012), .I2(n8752), .I3(n8751), .O(n8750) );
  ND2HHD U13058 ( .I1(n8209), .I2(n7809), .O(n12312) );
  ND2KHD U13059 ( .I1(n11713), .I2(n8992), .O(n13821) );
  AN3HHD U13060 ( .I1(n12564), .I2(n9625), .I3(n11503), .O(n10526) );
  INVNHD U13061 ( .I(n10206), .O(n8908) );
  NR2GHD U13062 ( .I1(n10907), .I2(n10906), .O(n12783) );
  BUFQHD U13063 ( .I(n9450), .O(n9449) );
  ND2DHD U13064 ( .I1(n6562), .I2(n12351), .O(n12352) );
  OAI12EHD U13065 ( .B1(n9389), .B2(n15416), .A1(n14606), .O(n6328) );
  NR2EHD U13066 ( .I1(n11452), .I2(n9689), .O(n9688) );
  OR3EHD U13067 ( .I1(n11312), .I2(n11452), .I3(n11193), .O(n10586) );
  ND2HHD U13068 ( .I1(n12790), .I2(n10825), .O(n12695) );
  NR2EHD U13069 ( .I1(n10447), .I2(n12695), .O(n10448) );
  OR3HHD U13070 ( .I1(n11433), .I2(n11452), .I3(n11432), .O(n11434) );
  AN3HHD U13071 ( .I1(n13822), .I2(n13821), .I3(n13820), .O(n13824) );
  NR2GHD U13072 ( .I1(n11046), .I2(n11045), .O(n12722) );
  ND3EHD U13073 ( .I1(n11703), .I2(n11702), .I3(_i_CLEFIA128_state_reg _1), .O(n11704) );
  MUX2HHD U13074 ( .A(n11698), .B(n11697), .S(_i_CLEFIA128_keyL _118), .O(n11703) );
  ND3CHD U13075 ( .I1(n12725), .I2(n11051), .I3(n11376), .O(n9702) );
  XOR2EHD U13076 ( .I1(DOUT_7), .I2(n6788), .O(n9970) );
  NR2EHD U13077 ( .I1(n11109), .I2(n11475), .O(n11114) );
  ND3EHD U13078 ( .I1(n11912), .I2(n11913), .I3(n13367), .O(n11926) );
  INVJHD U13079 ( .I(n9654), .O(n10244) );
  OR3HHD U13080 ( .I1(n12844), .I2(n12843), .I3(n12883), .O(n12845) );
  ND2HHD U13081 ( .I1(n8196), .I2(n8279), .O(n13680) );
  AN3EHD U13082 ( .I1(n7146), .I2(n10073), .I3(n11364), .O(n11047) );
  NR2GHD U13083 ( .I1(n11796), .I2(n11797), .O(n11798) );
  AN2HHD U13084 ( .I1(n8904), .I2(n11049), .O(n10074) );
  INVNHD U13085 ( .I(n8773), .O(n11049) );
  NR2EHD U13086 ( .I1(n11383), .I2(n11384), .O(n11385) );
  AN2HHD U13087 ( .I1(n12968), .I2(n12969), .O(n12973) );
  ND2HHD U13088 ( .I1(n11571), .I2(_i_CLEFIA128_state_reg _1), .O(n10189) );
  ND2KHD U13089 ( .I1(n9897), .I2(n9801), .O(n11491) );
  NR2GHD U13090 ( .I1(n12202), .I2(n12203), .O(n14074) );
  ND2HHD U13091 ( .I1(n13479), .I2(n13083), .O(n12202) );
  INVCHD U13092 ( .I(n10284), .O(n12784) );
  INVNHD U13093 ( .I(n9758), .O(n9800) );
  OR2KHD U13094 ( .I1(n8801), .I2(n11547), .O(n8759) );
  ND2HHD U13095 ( .I1(n9845), .I2(n11787), .O(n8818) );
  ND2KHD U13096 ( .I1(n12127), .I2(n11995), .O(n13629) );
  NR2IHD U13097 ( .I1(n11893), .I2(n12975), .O(n11892) );
  ND2KHD U13098 ( .I1(n12125), .I2(n12902), .O(n9772) );
  INVJHD U13099 ( .I(n8755), .O(n10160) );
  AN3EHD U13100 ( .I1(n13096), .I2(n14053), .I3(n8197), .O(n13092) );
  ND2KHD U13101 ( .I1(n9266), .I2(n9264), .O(n8763) );
  ND2KHD U13102 ( .I1(n7674), .I2(n8903), .O(n10484) );
  BUFEHD U13103 ( .I(n9127), .O(n9126) );
  ND2HHD U13104 ( .I1(n6959), .I2(n13550), .O(n9834) );
  XOR2EHD U13105 ( .I1(n14344), .I2(n8830), .O(n12138) );
  XOR2HHD U13106 ( .I1(n8764), .I2(n12828), .O(n10063) );
  ND2HHD U13107 ( .I1(n11673), .I2(_i_CLEFIA128_state_reg _1), .O(n11674) );
  INVCKGHD U13108 ( .I(n13419), .O(n11954) );
  AN3HHD U13109 ( .I1(n12582), .I2(n11358), .I3(n12559), .O(n12719) );
  NR2EHD U13110 ( .I1(n10937), .I2(n10744), .O(n9380) );
  XNR3EHD U13111 ( .I1(n8765), .I2(n14193), .I3(n14194), .O(n9755) );
  NR2IHD U13112 ( .I1(n8858), .I2(n11301), .O(n11464) );
  NR2EHD U13113 ( .I1(n12155), .I2(n13525), .O(n12156) );
  ND2HHD U13114 ( .I1(n9136), .I2(n11546), .O(n8770) );
  NR2GHD U13115 ( .I1(n13408), .I2(n12322), .O(n11941) );
  ND2HHD U13116 ( .I1(n11378), .I2(n9050), .O(n11379) );
  ND2KHD U13117 ( .I1(n11555), .I2(n12451), .O(n11168) );
  XNR2KHD U13118 ( .I1(n8772), .I2(n10162), .O(n12497) );
  INVGHD U13119 ( .I(n11318), .O(n10628) );
  ND3HHD U13120 ( .I1(n12742), .I2(n12564), .I3(n10485), .O(n11101) );
  BUFKHD U13121 ( .I(n10485), .O(n9625) );
  NR2EHD U13122 ( .I1(n12579), .I2(n11383), .O(n10530) );
  NR2EHD U13123 ( .I1(n9302), .I2(n9952), .O(n10831) );
  INVDHD U13124 ( .I(n12837), .O(n9468) );
  ND2HHD U13125 ( .I1(n9785), .I2(n9784), .O(n8774) );
  ND2KHD U13126 ( .I1(n9651), .I2(n7132), .O(n8792) );
  INVJHD U13127 ( .I(n6765), .O(n11417) );
  NR2GHD U13128 ( .I1(n11392), .I2(n11350), .O(n12571) );
  NR2CHD U13129 ( .I1(n9140), .I2(n9139), .O(n11184) );
  OR2KHD U13130 ( .I1(n7783), .I2(n10205), .O(n10206) );
  BUFQHD U13131 ( .I(n12004), .O(n13132) );
  ND2HHD U13132 ( .I1(n10959), .I2(n8979), .O(n10763) );
  NR2EHD U13133 ( .I1(n11532), .I2(n12470), .O(n11533) );
  ND2DHD U13134 ( .I1(n8938), .I2(n12794), .O(n10768) );
  OAI12EHD U13135 ( .B1(n12829), .B2(n10219), .A1(n8938), .O(n8920) );
  ND3EHD U13136 ( .I1(n11535), .I2(n11533), .I3(n11534), .O(n11538) );
  XNR2KHD U13137 ( .I1(n8788), .I2(n8793), .O(n14016) );
  ND2HHD U13138 ( .I1(n10037), .I2(n10145), .O(n9037) );
  BUFHHD U13139 ( .I(n9224), .O(n9222) );
  ND2HHD U13140 ( .I1(n8209), .I2(n7809), .O(n8779) );
  XNR2KHD U13141 ( .I1(n14489), .I2(n9958), .O(n12828) );
  INVGHD U13142 ( .I(n12309), .O(n11715) );
  OA13EHD U13143 ( .B1(n10725), .B2(n11137), .B3(n12508), .A1(n12506), .O(n10726) );
  NR2CHD U13144 ( .I1(n10586), .I2(n11537), .O(n8907) );
  ND2HHD U13145 ( .I1(n12454), .I2(n12469), .O(n10594) );
  ND2HHD U13146 ( .I1(n12730), .I2(n12564), .O(n11488) );
  ND2HHD U13147 ( .I1(n12687), .I2(n10448), .O(n10449) );
  ND3EHD U13148 ( .I1(n11808), .I2(n11809), .I3(n13533), .O(n11810) );
  INVJHD U13149 ( .I(n12836), .O(n12708) );
  ND2HHD U13150 ( .I1(n8797), .I2(_i_CLEFIA128_keyK _18), .O(n10562) );
  INVGHD U13151 ( .I(n9894), .O(n9351) );
  NR2CHD U13152 ( .I1(n9340), .I2(n9236), .O(n9339) );
  ND2DHD U13153 ( .I1(n9894), .I2(n10250), .O(n8783) );
  ND2HHD U13154 ( .I1(n7146), .I2(n7152), .O(n11118) );
  AN2HHD U13155 ( .I1(n10209), .I2(n12216), .O(n8784) );
  ND2HHD U13156 ( .I1(n10048), .I2(n10046), .O(n10045) );
  NR2GHD U13157 ( .I1(n11228), .I2(n10049), .O(n10048) );
  BUFQHD U13158 ( .I(n11976), .O(n12383) );
  OA112EHD U13159 ( .C1(n7166), .C2(n11222), .A1(n11221), .B1(n6803), .O(n8785) );
  ND3EHD U13160 ( .I1(n11781), .I2(n8341), .I3(n11780), .O(n11785) );
  NR2IHD U13161 ( .I1(n10631), .I2(n10630), .O(n11231) );
  ND2KHD U13162 ( .I1(n12092), .I2(n9235), .O(n9236) );
  ND2DHD U13163 ( .I1(n9035), .I2(n9038), .O(n8786) );
  ND2HHD U13164 ( .I1(n13512), .I2(n12302), .O(n13549) );
  ND3EHD U13165 ( .I1(n11145), .I2(n11147), .I3(n11146), .O(n11544) );
  ND2HHD U13166 ( .I1(n13102), .I2(n9556), .O(n11635) );
  BUFQHD U13167 ( .I(n11992), .O(n12129) );
  NR2EHD U13168 ( .I1(n13682), .I2(n13683), .O(n13685) );
  AN2HHD U13169 ( .I1(n9841), .I2(n8230), .O(n9651) );
  INVNHD U13170 ( .I(n8792), .O(n9801) );
  ND2HHD U13171 ( .I1(n13531), .I2(n13530), .O(n13553) );
  XOR2HHD U13172 ( .I1(n10140), .I2(n9912), .O(n8787) );
  ND2HHD U13173 ( .I1(n12402), .I2(n13613), .O(n12395) );
  ND3CHD U13174 ( .I1(n13144), .I2(n13143), .I3(n13187), .O(n13145) );
  ND2KHD U13175 ( .I1(n8225), .I2(n8889), .O(n9648) );
  ND2DHD U13176 ( .I1(n13844), .I2(n11814), .O(n9662) );
  ND3EHD U13177 ( .I1(n11348), .I2(n11347), .I3(n11346), .O(n11356) );
  ND2DHD U13178 ( .I1(n14053), .I2(n14082), .O(n9823) );
  ND2DHD U13179 ( .I1(n13088), .I2(n14082), .O(n13090) );
  ND2HHD U13180 ( .I1(n12327), .I2(n12351), .O(n12439) );
  AN2KHD U13181 ( .I1(n11300), .I2(n10628), .O(n12462) );
  ND2KHD U13182 ( .I1(n9626), .I2(n12484), .O(n11296) );
  AN3B1EHD U13183 ( .I1(n11491), .I2(n10073), .B1(n10074), .O(n11492) );
  BUFMHD U13184 ( .I(n13577), .O(n9747) );
  NR2CHD U13185 ( .I1(n10246), .I2(n11203), .O(n10288) );
  ND2HHD U13186 ( .I1(n7705), .I2(n11333), .O(n11034) );
  ND2HHD U13187 ( .I1(n9558), .I2(n13107), .O(n9718) );
  BUFMHD U13188 ( .I(n11416), .O(n9194) );
  ND2HHD U13189 ( .I1(n10850), .I2(n12609), .O(n12600) );
  BUFEHD U13190 ( .I(n14490), .O(n9757) );
  ND2HHD U13191 ( .I1(n11801), .I2(n7386), .O(n11802) );
  BUFQHD U13192 ( .I(n12363), .O(n9676) );
  XNR2KHD U13193 ( .I1(n14695), .I2(n14705), .O(n9867) );
  ND3CHD U13194 ( .I1(n13812), .I2(n13811), .I3(n13810), .O(n13813) );
  ND3CHD U13195 ( .I1(n11522), .I2(n11521), .I3(n11520), .O(n8880) );
  NR2EHD U13196 ( .I1(n12748), .I2(n11504), .O(n9103) );
  NR2EHD U13197 ( .I1(n11804), .I2(n11805), .O(n11809) );
  ND2HHD U13198 ( .I1(n12727), .I2(n12578), .O(n11471) );
  AN2HHD U13199 ( .I1(n13019), .I2(n13398), .O(n12331) );
  ND2DHD U13200 ( .I1(n12651), .I2(n12652), .O(n12654) );
  ND3EHD U13201 ( .I1(n11252), .I2(n11251), .I3(n9219), .O(n11258) );
  NR2GHD U13202 ( .I1(n8823), .I2(n11273), .O(n11314) );
  ND2DHD U13203 ( .I1(n12935), .I2(n12045), .O(n12277) );
  AN3EHD U13204 ( .I1(n14070), .I2(n10296), .I3(n9006), .O(n13055) );
  ND3CHD U13205 ( .I1(n13164), .I2(n13595), .I3(n9463), .O(n13166) );
  NR2GHD U13206 ( .I1(n13244), .I2(n11746), .O(n13491) );
  NR2EHD U13207 ( .I1(n12757), .I2(n9086), .O(n12570) );
  NR2IHD U13208 ( .I1(n10069), .I2(n10070), .O(n11484) );
  NR2GHD U13209 ( .I1(n11650), .I2(n8340), .O(n8795) );
  ND2HHD U13210 ( .I1(n13478), .I2(n9806), .O(n9569) );
  AN2EHD U13211 ( .I1(n13602), .I2(n12402), .O(n12293) );
  ND2DHD U13212 ( .I1(n7507), .I2(n10773), .O(n10775) );
  ND2KHD U13213 ( .I1(n8984), .I2(n8985), .O(n14167) );
  INVJHD U13214 ( .I(n7420), .O(n9991) );
  ND2DHD U13215 ( .I1(n10076), .I2(n15500), .O(n10001) );
  ND2KHD U13216 ( .I1(n9935), .I2(n9936), .O(n13911) );
  INVNHD U13217 ( .I(n9700), .O(n12561) );
  BUFQHD U13218 ( .I(n10480), .O(n11335) );
  NR2GHD U13219 ( .I1(n12108), .I2(n12107), .O(n12109) );
  ND3CHD U13220 ( .I1(n7118), .I2(n9806), .I3(n13096), .O(n11613) );
  ND2HHD U13221 ( .I1(n15134), .I2(n10292), .O(n13049) );
  ND2DHD U13222 ( .I1(n11292), .I2(n11541), .O(n11161) );
  NR2EHD U13223 ( .I1(n11000), .I2(n9968), .O(n9652) );
  BUFQHD U13224 ( .I(n10384), .O(n9659) );
  ND3CHD U13225 ( .I1(n9397), .I2(n11210), .I3(n11209), .O(n11211) );
  NR2CHD U13226 ( .I1(n11081), .I2(n11080), .O(n11082) );
  ND2HHD U13227 ( .I1(n12618), .I2(n11236), .O(n11059) );
  ND2HHD U13228 ( .I1(n11063), .I2(n12522), .O(n9261) );
  ND2HHD U13229 ( .I1(n7217), .I2(n9042), .O(n10776) );
  ND2HHD U13230 ( .I1(n12621), .I2(n9709), .O(n10789) );
  NR2IHD U13231 ( .I1(BSY), .I2(n14425), .O(n10928) );
  ND2HHD U13232 ( .I1(n13506), .I2(n8803), .O(n13679) );
  ND2KHD U13233 ( .I1(n10746), .I2(n7723), .O(n8812) );
  ND2CHD U13234 ( .I1(n12320), .I2(n8779), .O(n12170) );
  ND3EHD U13235 ( .I1(n6958), .I2(n8779), .I3(n13550), .O(n9815) );
  ND2HHD U13236 ( .I1(n8805), .I2(n13892), .O(n6104) );
  XNR2HHD U13237 ( .I1(DOUT_23), .I2(n9960), .O(n8806) );
  ND2HHD U13238 ( .I1(n8914), .I2(n12677), .O(n8810) );
  ND2HHD U13239 ( .I1(n10965), .I2(n8888), .O(n8811) );
  ND2HHD U13240 ( .I1(n8814), .I2(n10904), .O(n9871) );
  NR2IHD U13241 ( .I1(n7030), .I2(n8813), .O(n10904) );
  INVGHD U13242 ( .I(n8815), .O(n11799) );
  ND3EHD U13243 ( .I1(n12091), .I2(n13530), .I3(n13531), .O(n8817) );
  ND2KHD U13244 ( .I1(n12299), .I2(n12163), .O(n13682) );
  ND3EHD U13245 ( .I1(n8361), .I2(n8820), .I3(n11791), .O(n8819) );
  NR2BHD U13246 ( .I1(n8823), .I2(n12496), .O(n10716) );
  ND2KHD U13247 ( .I1(n11297), .I2(n11296), .O(n8823) );
  ND2CHD U13248 ( .I1(n8822), .I2(n10707), .O(n12495) );
  ND3EHD U13249 ( .I1(n11966), .I2(n8824), .I3(n8825), .O(n9984) );
  NR2EHD U13250 ( .I1(n8691), .I2(n9996), .O(n8827) );
  XOR2HHD U13251 ( .I1(_i_CLEFIA128_CON_T_x _10), .I2(DOUT_121), .O(n9996));
  OR3HHD U13252 ( .I1(n12188), .I2(n8828), .I3(n11749), .O(n11757) );
  OR3HHD U13253 ( .I1(n9696), .I2(n11771), .I3(n8828), .O(n11772) );
  NR2IHD U13254 ( .I1(n8833), .I2(n12216), .O(n11942) );
  NR2IHD U13255 ( .I1(n9051), .I2(n8833), .O(n12363) );
  ND2HHD U13256 ( .I1(n12410), .I2(n12361), .O(n13011) );
  ND2HHD U13257 ( .I1(n8260), .I2(n12092), .O(n9178) );
  ND2HHD U13258 ( .I1(n9631), .I2(n9006), .O(n9491) );
  ND2KHD U13259 ( .I1(n7034), .I2(n7907), .O(n9006) );
  INVDHD U13260 ( .I(n9006), .O(n13472) );
  ND2DHD U13261 ( .I1(n9006), .I2(n14072), .O(n13068) );
  ND2CHD U13262 ( .I1(n8431), .I2(n8235), .O(n10330) );
  OA13EHD U13263 ( .B1(n9179), .B2(n8847), .B3(n9400), .A1(n14067), .O(n9399));
  OA13EHD U13264 ( .B1(n11837), .B2(n11836), .B3(n8847), .A1(n14076), .O(n11838) );
  ND2HHD U13265 ( .I1(n14048), .I2(n11831), .O(n8847) );
  INVGHD U13266 ( .I(n8848), .O(n13511) );
  ND2HHD U13267 ( .I1(n13842), .I2(n9300), .O(n8848) );
  ND2KHD U13268 ( .I1(n10599), .I2(n11176), .O(n11440) );
  ND2HHD U13269 ( .I1(n7866), .I2(n8199), .O(n8853) );
  ND2HHD U13270 ( .I1(n8855), .I2(n15334), .O(n6156) );
  ND2HHD U13271 ( .I1(n13838), .I2(n13681), .O(n12143) );
  ND2KHD U13272 ( .I1(n9730), .I2(n9659), .O(n11070) );
  OR3HHD U13273 ( .I1(n10877), .I2(n12511), .I3(n10876), .O(n9257) );
  ND3EHD U13274 ( .I1(n9075), .I2(n9967), .I3(n9965), .O(n12815) );
  ND2KHD U13275 ( .I1(n10645), .I2(n9211), .O(n12627) );
  ND3EHD U13276 ( .I1(n10084), .I2(n11263), .I3(n11068), .O(n10869) );
  ND2KHD U13277 ( .I1(n9801), .I2(n9694), .O(n11411) );
  ND3EHD U13278 ( .I1(n12779), .I2(n9610), .I3(n12778), .O(n8864) );
  NR2CHD U13279 ( .I1(n10796), .I2(n9027), .O(n10797) );
  ND2KHD U13280 ( .I1(n8791), .I2(n10179), .O(n9423) );
  NR2CHD U13281 ( .I1(n11189), .I2(n11190), .O(n11197) );
  NR2GHD U13282 ( .I1(n10877), .I2(n11212), .O(n11220) );
  AN3HHD U13283 ( .I1(n7000), .I2(n7376), .I3(n7900), .O(n11526) );
  XNR2HHD U13284 ( .I1(DOUT_2), .I2(n9013), .O(n13924) );
  INVGHD U13285 ( .I(n12526), .O(n9656) );
  ND3EHD U13286 ( .I1(n10888), .I2(n10966), .I3(n12858), .O(n12675) );
  ND2HHD U13287 ( .I1(n9211), .I2(n12637), .O(n10796) );
  ND2HHD U13288 ( .I1(n11743), .I2(n14066), .O(n11658) );
  ND3EHD U13289 ( .I1(n14055), .I2(n13222), .I3(n14070), .O(n11751) );
  ND2DHD U13290 ( .I1(n14055), .I2(n7842), .O(n13104) );
  NR2GHD U13291 ( .I1(n10701), .I2(n11305), .O(n10702) );
  ND3EHD U13292 ( .I1(n12158), .I2(n12157), .I3(n12156), .O(n12167) );
  AN2HHD U13293 ( .I1(n13460), .I2(n13365), .O(n9438) );
  OR3HHD U13294 ( .I1(n10724), .I2(n9931), .I3(n10723), .O(n10725) );
  ND2HHD U13295 ( .I1(n11178), .I2(n9461), .O(n9931) );
  ND3EHD U13296 ( .I1(n12313), .I2(n11730), .I3(n13533), .O(n13657) );
  OA12HHD U13297 ( .B1(n10238), .B2(n12492), .A1(n12506), .O(n11559) );
  ND2HHD U13298 ( .I1(n9195), .I2(n8308), .O(n12492) );
  ND2KHD U13299 ( .I1(n9144), .I2(n11459), .O(n11448) );
  ND2KHD U13300 ( .I1(n14081), .I2(n9742), .O(n9367) );
  ND2KHD U13301 ( .I1(n10599), .I2(n12498), .O(n11530) );
  ND3CHD U13302 ( .I1(n11542), .I2(n11011), .I3(n11010), .O(n9919) );
  ND2KHD U13303 ( .I1(n9903), .I2(n9626), .O(n9443) );
  INVGHD U13304 ( .I(n12254), .O(n13032) );
  OA13EHD U13305 ( .B1(n13552), .B2(n13551), .B3(n13553), .A1(n8294), .O(n13554) );
  INVKHD U13306 ( .I(n9518), .O(n11648) );
  ND3EHD U13307 ( .I1(n10107), .I2(n12216), .I3(n10209), .O(n10291) );
  ND2HHD U13308 ( .I1(n10005), .I2(n13614), .O(n10006) );
  XOR2HHD U13309 ( .I1(n14138), .I2(n12815), .O(n9896) );
  ND2KHD U13310 ( .I1(n9730), .I2(n10874), .O(n12619) );
  AN3B1HHD U13311 ( .I1(n8197), .I2(n14070), .B1(n13473), .O(n12199) );
  OR3HHD U13312 ( .I1(n10861), .I2(n10833), .I3(n12648), .O(n8873) );
  XNR2KHD U13313 ( .I1(n10312), .I2(n8874), .O(n10325) );
  ND2HHD U13314 ( .I1(n8875), .I2(n15500), .O(n9079) );
  ND3EHD U13315 ( .I1(n11872), .I2(n11871), .I3(n11870), .O(n10110) );
  ND2KHD U13316 ( .I1(n6551), .I2(n8178), .O(n13659) );
  OR2KHD U13317 ( .I1(n12215), .I2(n9937), .O(n9706) );
  INVGHD U13318 ( .I(n12291), .O(n12292) );
  ND2HHD U13319 ( .I1(n8791), .I2(n7507), .O(n10645) );
  NR2IHD U13320 ( .I1(n12894), .I2(n8877), .O(n10079) );
  AN3HHD U13321 ( .I1(n12708), .I2(n10960), .I3(n10825), .O(n12792) );
  NR2IHD U13322 ( .I1(n9332), .I2(n10144), .O(n11677) );
  ND2KHD U13323 ( .I1(n11685), .I2(n9830), .O(n10144) );
  ND2HHD U13324 ( .I1(n8879), .I2(n12676), .O(n9975) );
  AN2HHD U13325 ( .I1(n12735), .I2(n10068), .O(n10066) );
  INVQHD U13326 ( .I(n8881), .O(n11995) );
  ND3EHD U13327 ( .I1(n12048), .I2(n6505), .I3(n13596), .O(n12049) );
  ND2KHD U13328 ( .I1(n8180), .I2(n11335), .O(n11358) );
  AN2HHD U13329 ( .I1(n8407), .I2(n11229), .O(n9584) );
  ND3EHD U13330 ( .I1(n9588), .I2(n12425), .I3(n12418), .O(n10104) );
  XNR2KHD U13331 ( .I1(n8378), .I2(n8885), .O(n10617) );
  INVNHD U13332 ( .I(_i_CLEFIA128_keyL _64), .O(n15408) );
  ND2HHD U13333 ( .I1(n11857), .I2(_i_CLEFIA128_keyL _107), .O(n8886) );
  OA13EHD U13334 ( .B1(n12509), .B2(n12507), .B3(n12508), .A1(n12506), .O(n9064) );
  ND3EHD U13335 ( .I1(n6997), .I2(n9708), .I3(n10022), .O(n10777) );
  NR2EHD U13336 ( .I1(n13146), .I2(n13145), .O(n13147) );
  ND2KHD U13337 ( .I1(n12423), .I2(n7058), .O(n12366) );
  ND3EHD U13338 ( .I1(n11210), .I2(n9618), .I3(n11204), .O(n9028) );
  NR2GHD U13339 ( .I1(n10789), .I2(n12600), .O(n11210) );
  ND3EHD U13340 ( .I1(n9726), .I2(n12951), .I3(n9093), .O(n12953) );
  ND3EHD U13341 ( .I1(n10029), .I2(n9412), .I3(n9410), .O(n9413) );
  INVGHD U13342 ( .I(n12186), .O(n9312) );
  OA13EHD U13343 ( .B1(n11543), .B2(n11545), .B3(n11544), .A1(n12491), .O(n11560) );
  ND2KHD U13344 ( .I1(n10179), .I2(n10318), .O(n10806) );
  ND2HHD U13345 ( .I1(n9604), .I2(n8178), .O(n12162) );
  ND3EHD U13346 ( .I1(n9030), .I2(n11777), .I3(n13804), .O(n11778) );
  ND2KHD U13347 ( .I1(n11713), .I2(n9435), .O(n12089) );
  NR2EHD U13348 ( .I1(n12229), .I2(n11894), .O(n11902) );
  OR3HHD U13349 ( .I1(n13446), .I2(n12412), .I3(n12413), .O(n12415) );
  ND2KHD U13350 ( .I1(n7034), .I2(n11834), .O(n9505) );
  ND3EHD U13351 ( .I1(n10740), .I2(n12690), .I3(n12677), .O(n10744) );
  NR2IHD U13352 ( .I1(n13115), .I2(n12117), .O(n12910) );
  AN2HHD U13353 ( .I1(n8893), .I2(n13835), .O(n10213) );
  ND3EHD U13354 ( .I1(n8894), .I2(n12315), .I3(n12316), .O(n8893) );
  ND3EHD U13355 ( .I1(n13135), .I2(n13134), .I3(n13182), .O(n13136) );
  NR2EHD U13356 ( .I1(n12256), .I2(n12255), .O(n12257) );
  OR3HHD U13357 ( .I1(n12937), .I2(n12938), .I3(n12936), .O(n12939) );
  INVCKGHD U13358 ( .I(n13184), .O(n13188) );
  XOR2HHD U13359 ( .I1(n9544), .I2(n13961), .O(n8898) );
  ND2KHD U13360 ( .I1(n9766), .I2(n10318), .O(n11262) );
  NR2GHD U13361 ( .I1(n9940), .I2(n9640), .O(n9939) );
  ND2HHD U13362 ( .I1(n8899), .I2(n8445), .O(n8987) );
  NR2CHD U13363 ( .I1(n11299), .I2(n9231), .O(n11304) );
  ND3EHD U13364 ( .I1(n12698), .I2(n12697), .I3(n12696), .O(n12699) );
  INVNHD U13365 ( .I(_i_CLEFIA128_keyL _16), .O(n15035) );
  XOR2HHD U13366 ( .I1(n14243), .I2(n6816), .O(n9956) );
  INVGHD U13367 ( .I(n11292), .O(n11141) );
  NR2IHD U13368 ( .I1(n10569), .I2(n11556), .O(n11523) );
  ND3EHD U13369 ( .I1(n6588), .I2(n12453), .I3(n12468), .O(n11136) );
  INVGHD U13370 ( .I(n10144), .O(n12173) );
  AN2HHD U13371 ( .I1(n12878), .I2(n12795), .O(n12798) );
  ND3EHD U13372 ( .I1(n10281), .I2(n8801), .I3(n10583), .O(n9681) );
  ND2HHD U13373 ( .I1(n11292), .I2(n12468), .O(n9196) );
  OA13EHD U13374 ( .B1(n11246), .B2(n11247), .B3(n12607), .A1(n6846), .O(n11269) );
  INVJHD U13375 ( .I(n9778), .O(n14766) );
  ND2KHD U13376 ( .I1(n10720), .I2(n10617), .O(n9110) );
  NR2EHD U13377 ( .I1(n13003), .I2(n13002), .O(n13009) );
  ND2HHD U13378 ( .I1(n10849), .I2(n12635), .O(n10663) );
  ND3EHD U13379 ( .I1(n8907), .I2(n8347), .I3(n8906), .O(n9647) );
  INVGHD U13380 ( .I(n8936), .O(n8935) );
  ND2KHD U13381 ( .I1(n8191), .I2(n8908), .O(n9003) );
  ND2KHD U13382 ( .I1(n10746), .I2(n8908), .O(n12692) );
  ND2KHD U13383 ( .I1(n10760), .I2(n8908), .O(n8914) );
  ND2HHD U13384 ( .I1(n10837), .I2(n8911), .O(n9601) );
  AN2HHD U13385 ( .I1(n12521), .I2(n12635), .O(n8911) );
  INVCHD U13386 ( .I(n8914), .O(n8912) );
  BUFQHD U13387 ( .I(n9384), .O(n8916) );
  INVCKGHD U13388 ( .I(n9008), .O(n8922) );
  ND2HHD U13389 ( .I1(n9003), .I2(n12673), .O(n12665) );
  ND2HHD U13390 ( .I1(n9003), .I2(n10966), .O(n10750) );
  ND3EHD U13391 ( .I1(n8399), .I2(n8925), .I3(n8924), .O(n12787) );
  INVCKGHD U13392 ( .I(n12675), .O(n8924) );
  ND2HHD U13393 ( .I1(n8928), .I2(n8929), .O(n8927) );
  AN2HHD U13394 ( .I1(n8932), .I2(n8933), .O(n8931) );
  ND2HHD U13395 ( .I1(n9991), .I2(n12713), .O(n8932) );
  ND2HHD U13396 ( .I1(n9993), .I2(n10088), .O(n8933) );
  XOR2EHD U13397 ( .I1(n8793), .I2(n9255), .O(n13923) );
  ND3EHD U13398 ( .I1(n8940), .I2(n8943), .I3(n8941), .O(n8939) );
  OR2HHD U13399 ( .I1(n10946), .I2(n10943), .O(n8954) );
  ND2HHD U13400 ( .I1(n8956), .I2(n10970), .O(n8955) );
  NR2GHD U13401 ( .I1(n8959), .I2(n8958), .O(n10740) );
  ND2KHD U13402 ( .I1(n8961), .I2(n8960), .O(n10825) );
  ND2HHD U13403 ( .I1(n8962), .I2(n12690), .O(n9454) );
  ND2HHD U13404 ( .I1(n10990), .I2(n8976), .O(n11156) );
  ND2CHD U13405 ( .I1(n12469), .I2(n8976), .O(n11442) );
  ND2HHD U13406 ( .I1(n9531), .I2(n8976), .O(n9953) );
  ND2KHD U13407 ( .I1(n10973), .I2(n11274), .O(n8976) );
  NR2GHD U13408 ( .I1(n8978), .I2(n10812), .O(n10813) );
  ND2CHD U13409 ( .I1(n9669), .I2(n8979), .O(n10829) );
  ND2KHD U13410 ( .I1(n9581), .I2(n9383), .O(n10965) );
  ND2KHD U13411 ( .I1(n10124), .I2(n10738), .O(n12790) );
  XOR2HHD U13412 ( .I1(n10232), .I2(n8981), .O(n10230) );
  INVQHD U13413 ( .I(_i_CLEFIA128_keyL _101), .O(n8982) );
  OR2EHD U13414 ( .I1(n8797), .I2(n8982), .O(n11970) );
  ND2KHD U13415 ( .I1(n10452), .I2(n10939), .O(n12876) );
  ND3EHD U13416 ( .I1(n6993), .I2(n8344), .I3(n8983), .O(n12510) );
  XNR3EHD U13417 ( .I1(n8988), .I2(n10180), .I3(n14367), .O(n9078) );
  ND2HHD U13418 ( .I1(n8989), .I2(n13431), .O(n9249) );
  ND3EHD U13419 ( .I1(n9254), .I2(n9253), .I3(n9250), .O(n8989) );
  ND2DHD U13420 ( .I1(n12291), .I2(n12901), .O(n13144) );
  ND2KHD U13421 ( .I1(n12411), .I2(n7114), .O(n12989) );
  ND2KHD U13422 ( .I1(n11906), .I2(n9449), .O(n13383) );
  ND3EHD U13423 ( .I1(n10009), .I2(n10222), .I3(n13212), .O(n13169) );
  ND3EHD U13424 ( .I1(n12999), .I2(n13022), .I3(n13021), .O(n13461) );
  ND2HHD U13425 ( .I1(n9167), .I2(n9170), .O(n8994) );
  ND2KHD U13426 ( .I1(n11766), .I2(n9183), .O(n14055) );
  ND2HHD U13427 ( .I1(n13399), .I2(n13021), .O(n12360) );
  ND2KHD U13428 ( .I1(n9626), .I2(n12498), .O(n11546) );
  BUFNHD U13429 ( .I(n9455), .O(n9184) );
  ND2HHD U13430 ( .I1(n9009), .I2(n9440), .O(n6107) );
  NR2CHD U13431 ( .I1(n12695), .I2(n12807), .O(n12696) );
  BUFNHD U13432 ( .I(n10007), .O(n10005) );
  NR2EHD U13433 ( .I1(n9155), .I2(n10261), .O(n9154) );
  ND2HHD U13434 ( .I1(n8995), .I2(n9567), .O(n10140) );
  ND3EHD U13435 ( .I1(n9111), .I2(n7003), .I3(n7002), .O(n11537) );
  ND2HHD U13436 ( .I1(n9443), .I2(n12454), .O(n10572) );
  OA12HHD U13437 ( .B1(n9827), .B2(n9828), .A1(n13835), .O(n9826) );
  BUFMHD U13438 ( .I(n9237), .O(n9072) );
  NR2IHD U13439 ( .I1(n11066), .I2(n10362), .O(n11232) );
  ND2KHD U13440 ( .I1(n13640), .I2(n13641), .O(n14028) );
  NR2IHD U13441 ( .I1(n11126), .I2(n9751), .O(n10215) );
  OA12HHD U13442 ( .B1(n11387), .B2(n11388), .A1(n11500), .O(n11389) );
  ND3EHD U13443 ( .I1(n10783), .I2(n10862), .I3(n10851), .O(n11259) );
  ND3EHD U13444 ( .I1(n13866), .I2(n13868), .I3(n13867), .O(n6166) );
  ND2HHD U13445 ( .I1(n12616), .I2(n12615), .O(n12649) );
  INVGHD U13446 ( .I(n10005), .O(n13574) );
  ND2KHD U13447 ( .I1(n12900), .I2(n9580), .O(n9832) );
  ND2KHD U13448 ( .I1(n9684), .I2(n10760), .O(n12689) );
  XNR2HHD U13449 ( .I1(n11695), .I2(n11694), .O(n11736) );
  XNR2HHD U13450 ( .I1(n11705), .I2(n11704), .O(n11737) );
  ND3EHD U13451 ( .I1(n10542), .I2(n9716), .I3(n10543), .O(n9010) );
  AN2HHD U13452 ( .I1(n11727), .I2(n11737), .O(n13817) );
  NR2EHD U13453 ( .I1(n12404), .I2(n12403), .O(n12405) );
  OA13EHD U13454 ( .B1(n11106), .B2(n11107), .B3(n9534), .A1(n12591), .O(n9751) );
  ND2HHD U13455 ( .I1(n13789), .I2(n13788), .O(n6111) );
  ND2KHD U13456 ( .I1(n7621), .I2(n12484), .O(n12478) );
  BUFQHD U13457 ( .I(n11943), .O(n9430) );
  ND2HHD U13458 ( .I1(n9072), .I2(n9136), .O(n11193) );
  ND2KHD U13459 ( .I1(n6872), .I2(n12145), .O(n12299) );
  ND2KHD U13460 ( .I1(n6909), .I2(n8214), .O(n13000) );
  AN3HHD U13461 ( .I1(n9627), .I2(n12464), .I3(n12486), .O(n10596) );
  OAI112BHD U13462 ( .C1(n10096), .C2(n14378), .A1(n9018), .B1(n14387), .O(n6138) );
  BUFKHD U13463 ( .I(n12480), .O(n9047) );
  ND2KHD U13464 ( .I1(n12456), .I2(n11192), .O(n11280) );
  NR2EHD U13465 ( .I1(n12642), .I2(n12641), .O(n12643) );
  ND3EHD U13466 ( .I1(n12645), .I2(n12643), .I3(n12644), .O(n12647) );
  XOR2HHD U13467 ( .I1(n6808), .I2(n7256), .O(n9023) );
  ND2HHD U13468 ( .I1(n12166), .I2(n12165), .O(n13663) );
  NR2CHD U13469 ( .I1(n12326), .I2(n12325), .O(n12332) );
  AN2HHD U13470 ( .I1(n13396), .I2(n9398), .O(n13457) );
  BUFIHD U13471 ( .I(n11530), .O(n9053) );
  OA12HHD U13472 ( .B1(n11906), .B2(n12363), .A1(n7032), .O(n11957) );
  INVJHD U13473 ( .I(n9028), .O(n11078) );
  ND2HHD U13474 ( .I1(n14044), .I2(n11646), .O(n12211) );
  ND2HHD U13475 ( .I1(n12812), .I2(n12810), .O(n9347) );
  NR2EHD U13476 ( .I1(n12954), .I2(n12953), .O(n12959) );
  OR3HHD U13477 ( .I1(n9234), .I2(n9233), .I3(n9563), .O(n12232) );
  BUFEHD U13478 ( .I(n11843), .O(n9029) );
  NR2EHD U13479 ( .I1(n11734), .I2(n13830), .O(n11735) );
  BUFKHD U13480 ( .I(n12309), .O(n9030) );
  INVMHD U13481 ( .I(n9681), .O(n10600) );
  ND3CHD U13482 ( .I1(n12478), .I2(n12464), .I3(n9135), .O(n12465) );
  ND2HHD U13483 ( .I1(n11117), .I2(n10485), .O(n11092) );
  OA12HHD U13484 ( .B1(n10175), .B2(n11329), .A1(n12752), .O(n9033) );
  NR2GHD U13485 ( .I1(n13150), .I2(n13151), .O(n13155) );
  ND2HHD U13486 ( .I1(n9694), .I2(n11336), .O(n11482) );
  ND2KHD U13487 ( .I1(n10644), .I2(n7864), .O(n11079) );
  NR2EHD U13488 ( .I1(n8993), .I2(n11654), .O(n11655) );
  OA22HHD U13489 ( .A1(n9570), .A2(n11659), .B1(n11637), .B2(n13075), .O(n9035) );
  ND2HHD U13490 ( .I1(n13078), .I2(n13077), .O(n13079) );
  ND3EHD U13491 ( .I1(n12999), .I2(n12955), .I3(n12410), .O(n12334) );
  ND2KHD U13492 ( .I1(n7038), .I2(n9430), .O(n12999) );
  ND3EHD U13493 ( .I1(n9039), .I2(n9727), .I3(n12136), .O(n9040) );
  AN2HHD U13494 ( .I1(n9218), .I2(n11459), .O(n11460) );
  ND2KHD U13495 ( .I1(n9044), .I2(n9043), .O(n12298) );
  XNR2HHD U13496 ( .I1(DOUT_12), .I2(n14137), .O(n12886) );
  ND2KHD U13497 ( .I1(n11818), .I2(n11834), .O(n13098) );
  ND2HHD U13498 ( .I1(n13948), .I2(n13947), .O(n6142) );
  NR2IHD U13499 ( .I1(n11406), .I2(n11470), .O(n12735) );
  OR3EHD U13500 ( .I1(n12461), .I2(n9388), .I3(n12460), .O(n10272) );
  AN4EHD U13501 ( .I1(n13613), .I2(n13207), .I3(n13573), .I4(n13629), .O(n11994) );
  BUFKHD U13502 ( .I(n10208), .O(n9051) );
  BUFQHD U13503 ( .I(n14059), .O(n9597) );
  ND2KHD U13504 ( .I1(n9898), .I2(n7039), .O(n12553) );
  ND2KHD U13505 ( .I1(n12829), .I2(n9559), .O(n12688) );
  INVDHD U13506 ( .I(n11262), .O(n9055) );
  ND2HHD U13507 ( .I1(n9058), .I2(n9057), .O(n10092) );
  NR2GHD U13508 ( .I1(n10093), .I2(n13434), .O(n9057) );
  ND3EHD U13509 ( .I1(n10846), .I2(n6921), .I3(n10845), .O(n10852) );
  NR2GHD U13510 ( .I1(n9059), .I2(n9060), .O(n10438) );
  AN3HHD U13511 ( .I1(n10435), .I2(n7102), .I3(n9061), .O(n9060) );
  INVGHD U13512 ( .I(n13507), .O(n9177) );
  OR2EHD U13513 ( .I1(n6813), .I2(n12606), .O(n9063) );
  ND3EHD U13514 ( .I1(n10395), .I2(n10396), .I3(_i_CLEFIA128_state_reg _1), .O(n10397) );
  AN3HHD U13515 ( .I1(n10198), .I2(n8800), .I3(n11647), .O(n9455) );
  ND3EHD U13516 ( .I1(n9135), .I2(n11430), .I3(n9443), .O(n12503) );
  ND3EHD U13517 ( .I1(n12772), .I2(n6956), .I3(n12771), .O(n12773) );
  ND2DHD U13518 ( .I1(n10080), .I2(n12402), .O(n12097) );
  OR3HHD U13519 ( .I1(n13665), .I2(n13663), .I3(n13664), .O(n13667) );
  ND2HHD U13520 ( .I1(n13541), .I2(n12306), .O(n12308) );
  AN3HHD U13521 ( .I1(n9065), .I2(n10097), .I3(n10101), .O(n9686) );
  OAI12CHD U13522 ( .B1(n9889), .B2(n13437), .A1(n13458), .O(n9065) );
  ND2KHD U13523 ( .I1(n10178), .I2(n7864), .O(n10855) );
  ND2HHD U13524 ( .I1(n8416), .I2(n14048), .O(n9354) );
  INVDHD U13525 ( .I(n9125), .O(n9265) );
  AN2KHD U13526 ( .I1(n13577), .I2(n13199), .O(n12928) );
  ND3EHD U13527 ( .I1(n13076), .I2(n11841), .I3(n11842), .O(n12183) );
  AN2HHD U13528 ( .I1(n6932), .I2(n6935), .O(n13474) );
  XOR2HHD U13529 ( .I1(n14490), .I2(n13951), .O(n9959) );
  ND2HHD U13530 ( .I1(n13727), .I2(n13726), .O(n6126) );
  XOR3EHD U13531 ( .I1(n13716), .I2(n9550), .I3(n13753), .O(n15200) );
  INVMHD U13532 ( .I(n9645), .O(n13386) );
  ND2HHD U13533 ( .I1(n13066), .I2(n9742), .O(n13490) );
  INVQHD U13534 ( .I(_i_CLEFIA128_keyL _98), .O(n15120) );
  INVKHD U13535 ( .I(n9675), .O(n13430) );
  AN2HHD U13536 ( .I1(n13153), .I2(n13175), .O(n12406) );
  NR2EHD U13537 ( .I1(n10482), .I2(n11495), .O(n11100) );
  NR2GHD U13538 ( .I1(n15513), .I2(n9389), .O(n14347) );
  OR2EHD U13539 ( .I1(n12404), .I2(n12295), .O(n9070) );
  OR2HHD U13540 ( .I1(n13105), .I2(n13104), .O(n9485) );
  INVGHD U13541 ( .I(n12721), .O(n12723) );
  INVGHD U13542 ( .I(n11488), .O(n11489) );
  AN2HHD U13543 ( .I1(n12877), .I2(n12692), .O(n10421) );
  ND2HHD U13544 ( .I1(_i_CLEFIA128_keyK _4), .I2(_i_CLEFIA128_keyL _4), .O(n10458) );
  ND2KHD U13545 ( .I1(n12423), .I2(n9917), .O(n9679) );
  ND2KHD U13546 ( .I1(n11681), .I2(n7035), .O(n13804) );
  ND2KHD U13547 ( .I1(_i_CLEFIA128_keyK _108), .I2(n8797), .O(n11862) );
  XNR2HHD U13548 ( .I1(DOUT_13), .I2(n9761), .O(n14104) );
  ND2KHD U13549 ( .I1(n8797), .I2(_i_CLEFIA128_keyK _82), .O(n10563) );
  ND2HHD U13550 ( .I1(n9077), .I2(n9079), .O(n6210) );
  OR3HHD U13551 ( .I1(n9507), .I2(n11621), .I3(n11622), .O(n11623) );
  ND3EHD U13552 ( .I1(n8353), .I2(n9080), .I3(n9281), .O(n9280) );
  NR2EHD U13553 ( .I1(n9081), .I2(n9282), .O(n9080) );
  INVDHD U13554 ( .I(n9493), .O(n13100) );
  ND2HHD U13555 ( .I1(n15481), .I2(n15500), .O(n15485) );
  OAI112BHD U13556 ( .C1(n7831), .C2(n13691), .A1(n9082), .B1(n13698), .O(n6128) );
  ND2HHD U13557 ( .I1(n7831), .I2(n8268), .O(n9082) );
  ND2KHD U13558 ( .I1(n9807), .I2(n8196), .O(n13512) );
  ND2KHD U13559 ( .I1(n8771), .I2(n9549), .O(n13671) );
  INVKHD U13560 ( .I(n9085), .O(n12425) );
  ND2HHD U13561 ( .I1(n13399), .I2(n13028), .O(n9085) );
  ND2KHD U13562 ( .I1(n9699), .I2(n13132), .O(n13195) );
  OR3HHD U13563 ( .I1(n13587), .I2(n9629), .I3(n12926), .O(n12927) );
  ND2HHD U13564 ( .I1(n11335), .I2(n9694), .O(n10534) );
  ND2KHD U13565 ( .I1(n7254), .I2(n8178), .O(n13805) );
  AN2HHD U13566 ( .I1(n11646), .I2(n8254), .O(n12198) );
  ND3EHD U13567 ( .I1(n10722), .I2(n11464), .I3(n9088), .O(n12508) );
  OA12HHD U13568 ( .B1(n14621), .B2(n11129), .A1(n14196), .O(n14197) );
  ND3EHD U13569 ( .I1(n9090), .I2(n9221), .I3(n13370), .O(n12416) );
  XOR2HHD U13570 ( .I1(n14108), .I2(n7935), .O(n14006) );
  ND2HHD U13571 ( .I1(n13417), .I2(n13418), .O(n14108) );
  OAI22CHD U13572 ( .A1(n12291), .A2(n12900), .B1(n12383), .B2(n12127), .O(n12128) );
  NR2EHD U13573 ( .I1(n13385), .I2(n13384), .O(n13387) );
  ND3EHD U13574 ( .I1(n12620), .I2(n10673), .I3(n10850), .O(n11085) );
  ND3EHD U13575 ( .I1(n10706), .I2(n11307), .I3(n10707), .O(n11013) );
  ND2KHD U13576 ( .I1(n12900), .I2(n13132), .O(n13577) );
  OR3HHD U13577 ( .I1(n9525), .I2(n13828), .I3(n11720), .O(n9827) );
  OR3HHD U13578 ( .I1(n11712), .I2(n11710), .I3(n11711), .O(n13828) );
  ND2KHD U13579 ( .I1(n12030), .I2(n9580), .O(n10007) );
  AN3HHD U13580 ( .I1(n12877), .I2(n10961), .I3(n10962), .O(n10963) );
  ND2KHD U13581 ( .I1(n9684), .I2(n9383), .O(n12668) );
  INVMHD U13582 ( .I(_i_CLEFIA128_keyK _116), .O(n14377) );
  ND2HHD U13583 ( .I1(n12688), .I2(n10768), .O(n10769) );
  ND3EHD U13584 ( .I1(n10105), .I2(n10102), .I3(n12236), .O(n9096) );
  ND2KHD U13585 ( .I1(n11906), .I2(n9430), .O(n13401) );
  NR2GHD U13586 ( .I1(n11952), .I2(n9097), .O(n12254) );
  NR2IHD U13587 ( .I1(n11991), .I2(n6881), .O(n11976) );
  ND2KHD U13588 ( .I1(n13419), .I2(n13022), .O(n9645) );
  ND2KHD U13589 ( .I1(n14056), .I2(n9605), .O(n13243) );
  ND3EHD U13590 ( .I1(n9589), .I2(n8876), .I3(n8320), .O(n11939) );
  AN2HHD U13591 ( .I1(n9593), .I2(n12448), .O(n12452) );
  AN2HHD U13592 ( .I1(n13541), .I2(n13681), .O(n9235) );
  ND2KHD U13593 ( .I1(n11274), .I2(n12498), .O(n12449) );
  ND2HHD U13594 ( .I1(n9190), .I2(n12677), .O(n10766) );
  OA112HHD U13595 ( .C1(n11325), .C2(n11324), .A1(n12747), .B1(n12559), .O(n11326) );
  ND2KHD U13596 ( .I1(n9103), .I2(n6941), .O(n10073) );
  ND2DHD U13597 ( .I1(n12915), .I2(n8185), .O(n13164) );
  NR2GHD U13598 ( .I1(n12940), .I2(n12939), .O(n12943) );
  NR2IHD U13599 ( .I1(n11615), .I2(n11609), .O(n13097) );
  NR2EHD U13600 ( .I1(n11732), .I2(n11733), .O(n12149) );
  NR2EHD U13601 ( .I1(n9138), .I2(n9143), .O(n9137) );
  OR2KHD U13602 ( .I1(n8858), .I2(n9292), .O(n9291) );
  ND2KHD U13603 ( .I1(n10179), .I2(n9730), .O(n12521) );
  NR2CHD U13604 ( .I1(n9953), .I2(n10616), .O(n10623) );
  OAI112BHD U13605 ( .C1(n15449), .C2(n14032), .A1(n9106), .B1(n14039), .O(n6144) );
  ND2HHD U13606 ( .I1(n15449), .I2(n8269), .O(n9106) );
  ND3CHD U13607 ( .I1(n12191), .I2(n9806), .I3(n12192), .O(n12193) );
  ND3EHD U13608 ( .I1(n11718), .I2(n13677), .I3(n11719), .O(n11720) );
  ND2HHD U13609 ( .I1(n9108), .I2(n9107), .O(n6219) );
  NR2GHD U13610 ( .I1(n15513), .I2(n10008), .O(n9109) );
  BUFQHD U13611 ( .I(n11997), .O(n12902) );
  ND3EHD U13612 ( .I1(n10239), .I2(n11557), .I3(n11558), .O(n10238) );
  AN2HHD U13613 ( .I1(n10295), .I2(n12431), .O(n12432) );
  ND3EHD U13614 ( .I1(n9247), .I2(n9248), .I3(n12992), .O(n13039) );
  OR3HHD U13615 ( .I1(n9876), .I2(n12378), .I3(n13152), .O(n12379) );
  ND2HHD U13616 ( .I1(n12276), .I2(n12920), .O(n13152) );
  OA13EHD U13617 ( .B1(n13149), .B2(n13170), .B3(n9728), .A1(n13585), .O(n13159) );
  OR3HHD U13618 ( .I1(n13462), .I2(n13461), .I3(n13463), .O(n13464) );
  ND2HHD U13619 ( .I1(n9627), .I2(n9116), .O(n11160) );
  ND2CHD U13620 ( .I1(n9116), .I2(n9072), .O(n10616) );
  ND2CHD U13621 ( .I1(n11295), .I2(n9116), .O(n10977) );
  ND2HHD U13622 ( .I1(n11187), .I2(n9115), .O(n11190) );
  AN2CHD U13623 ( .I1(n9116), .I2(n11553), .O(n9115) );
  ND2KHD U13624 ( .I1(n7621), .I2(n11176), .O(n9116) );
  AN3HHD U13625 ( .I1(n12362), .I2(n8320), .I3(n13430), .O(n9117) );
  ND2KHD U13626 ( .I1(n8209), .I2(n9435), .O(n9759) );
  ND2KHD U13627 ( .I1(n9118), .I2(n13383), .O(n12359) );
  ND2KHD U13628 ( .I1(n6909), .I2(n9642), .O(n9118) );
  INVCKGHD U13629 ( .I(n9118), .O(n13016) );
  ND2CHD U13630 ( .I1(n9119), .I2(n9239), .O(n12246) );
  ND2KHD U13631 ( .I1(n11906), .I2(n7830), .O(n9119) );
  ND2HHD U13632 ( .I1(n9119), .I2(n12419), .O(n12420) );
  ND2HHD U13633 ( .I1(n13013), .I2(n9121), .O(n9120) );
  OR3HHD U13634 ( .I1(n11957), .I2(n11956), .I3(n9387), .O(n9973) );
  OR3HHD U13635 ( .I1(n13016), .I2(n13449), .I3(n13015), .O(n9124) );
  ND3EHD U13636 ( .I1(n13460), .I2(n13447), .I3(n13365), .O(n12441) );
  ND3EHD U13637 ( .I1(n6979), .I2(n6607), .I3(n9026), .O(n12227) );
  ND2CHD U13638 ( .I1(n13590), .I2(n9126), .O(n12135) );
  ND2KHD U13639 ( .I1(n10095), .I2(n12129), .O(n9127) );
  ND2HHD U13640 ( .I1(n8216), .I2(n6873), .O(n9128) );
  ND2CHD U13641 ( .I1(n9129), .I2(n6553), .O(n11285) );
  INVLHD U13642 ( .I(_i_CLEFIA128_keyL _84), .O(n15089) );
  OAI12CHD U13643 ( .B1(n10096), .B2(n15416), .A1(n14668), .O(n6265) );
  ND2HHD U13644 ( .I1(n9136), .I2(n11553), .O(n11433) );
  ND2HHD U13645 ( .I1(n11552), .I2(n9136), .O(n11283) );
  ND2KHD U13646 ( .I1(n9964), .I2(n12498), .O(n9136) );
  ND2HHD U13647 ( .I1(n9137), .I2(n11307), .O(n11135) );
  ND3EHD U13648 ( .I1(n9297), .I2(n12464), .I3(n12450), .O(n9296) );
  ND2HHD U13649 ( .I1(n9141), .I2(n13740), .O(n6110) );
  XOR2HHD U13650 ( .I1(n13730), .I2(n9142), .O(n14573) );
  XOR2HHD U13651 ( .I1(n13731), .I2(n9550), .O(n9142) );
  ND2CHD U13652 ( .I1(n9593), .I2(n9144), .O(n10698) );
  ND2KHD U13653 ( .I1(n12498), .I2(n9800), .O(n9144) );
  ND2HHD U13654 ( .I1(n9145), .I2(n9709), .O(n10356) );
  ND2KHD U13655 ( .I1(n7217), .I2(n10874), .O(n9145) );
  ND2DHD U13656 ( .I1(n9151), .I2(n7043), .O(n9147) );
  OAI112BHD U13657 ( .C1(n9151), .C2(n8388), .A1(n9148), .B1(n13960), .O(n6113) );
  ND3EHD U13658 ( .I1(n15454), .I2(n9150), .I3(n15453), .O(n6204) );
  ND2HHD U13659 ( .I1(n9160), .I2(n9158), .O(n14141) );
  ND3EHD U13660 ( .I1(n9162), .I2(n9360), .I3(n9159), .O(n9158) );
  AN2HHD U13661 ( .I1(n11458), .I2(n12491), .O(n9161) );
  OA13EHD U13662 ( .B1(n11428), .B2(n12475), .B3(n11427), .A1(n12474), .O(n9163) );
  OA12HHD U13663 ( .B1(n12463), .B2(n9798), .A1(n12506), .O(n9164) );
  ND2CHD U13664 ( .I1(n13182), .I2(n12935), .O(n12937) );
  OR2EHD U13665 ( .I1(n9166), .I2(n13171), .O(n13174) );
  ND2CHD U13666 ( .I1(n12123), .I2(n13182), .O(n9166) );
  NR2GHD U13667 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(n9174), .O(n9168) );
  NR2EHD U13668 ( .I1(n9175), .I2(n9720), .O(n9170) );
  XNR2KHD U13669 ( .I1(_i_CLEFIA128_keyL _115), .I2(n11667), .O(n9174) );
  AN2HHD U13670 ( .I1(n9177), .I2(n11730), .O(n12315) );
  OR3HHD U13671 ( .I1(n14058), .I2(n9180), .I3(n14064), .O(n9179) );
  ND3EHD U13672 ( .I1(n9181), .I2(n14081), .I3(n14063), .O(n9180) );
  NR2GHD U13673 ( .I1(n11829), .I2(n11830), .O(n14048) );
  NR2GHD U13674 ( .I1(n9920), .I2(n9921), .O(n11831) );
  BUFNHD U13675 ( .I(n9422), .O(n9183) );
  AN2HHD U13676 ( .I1(n9185), .I2(n14063), .O(n13482) );
  ND2HHD U13677 ( .I1(n9190), .I2(n12688), .O(n12800) );
  ND2HHD U13678 ( .I1(n12832), .I2(n9190), .O(n12670) );
  ND2CHD U13679 ( .I1(n10960), .I2(n9190), .O(n10894) );
  ND2KHD U13680 ( .I1(n10874), .I2(n10178), .O(n9191) );
  ND3EHD U13681 ( .I1(n10783), .I2(n11225), .I3(n9191), .O(n10662) );
  OR2B1CHD U13682 ( .I1(n10836), .B1(n12598), .O(n12599) );
  ND2HHD U13683 ( .I1(n6841), .I2(n11262), .O(n12614) );
  XOR2HHD U13684 ( .I1(_i_CLEFIA128_keyL _83), .I2(n9193), .O(n10550) );
  ND2KHD U13685 ( .I1(n9904), .I2(n9905), .O(n9961) );
  OR3HHD U13686 ( .I1(n9197), .I2(n11715), .I3(n11714), .O(n9525) );
  OA13EHD U13687 ( .B1(n9198), .B2(n13544), .B3(n13545), .A1(n13826), .O(n13555) );
  OA13EHD U13688 ( .B1(n13534), .B2(n9198), .B3(n13553), .A1(n13817), .O(n13535) );
  ND2KHD U13689 ( .I1(n9199), .I2(n13533), .O(n9434) );
  ND2CHD U13690 ( .I1(n6766), .I2(n10973), .O(n10974) );
  ND2KHD U13691 ( .I1(n10973), .I2(n6873), .O(n12501) );
  XNR2KHD U13692 ( .I1(n10551), .I2(n9202), .O(n10587) );
  AN2HHD U13693 ( .I1(n9205), .I2(_i_CLEFIA128_state_reg _1), .O(n9204) );
  ND2KHD U13694 ( .I1(n7161), .I2(n6882), .O(n9211) );
  NR2CHD U13695 ( .I1(n9213), .I2(n9212), .O(n13433) );
  ND2HHD U13696 ( .I1(n9216), .I2(n9311), .O(n10210) );
  ND2CHD U13697 ( .I1(n12253), .I2(n9216), .O(n13376) );
  ND3CHD U13698 ( .I1(n12986), .I2(n12987), .I3(n9216), .O(n12993) );
  XNR2KHD U13699 ( .I1(n10555), .I2(n10554), .O(n10281) );
  ND2KHD U13700 ( .I1(n11530), .I2(n9218), .O(n12496) );
  AN2HHD U13701 ( .I1(n12533), .I2(n9219), .O(n12534) );
  OA12HHD U13702 ( .B1(n9220), .B2(n12074), .A1(n13826), .O(n9824) );
  NR2IHD U13703 ( .I1(n9706), .I2(n9707), .O(n9221) );
  ND2KHD U13704 ( .I1(n9224), .I2(n11554), .O(n11305) );
  ND2DHD U13705 ( .I1(n9443), .I2(n9224), .O(n9223) );
  ND2CHD U13706 ( .I1(n9224), .I2(n12469), .O(n11009) );
  ND2KHD U13707 ( .I1(n9626), .I2(n10600), .O(n9224) );
  INVCHD U13708 ( .I(n12423), .O(n9225) );
  XOR2HHD U13709 ( .I1(DOUT_95), .I2(n9923), .O(n9710) );
  ND2HHD U13710 ( .I1(n11758), .I2(n8348), .O(n11753) );
  ND2HHD U13711 ( .I1(n9229), .I2(n7001), .O(n9555) );
  ND3EHD U13712 ( .I1(n9462), .I2(n9185), .I3(n11649), .O(n11650) );
  ND3CHD U13713 ( .I1(n9006), .I2(n13217), .I3(n9462), .O(n9921) );
  ND2KHD U13714 ( .I1(n7292), .I2(n8078), .O(n9462) );
  OR3HHD U13715 ( .I1(n11168), .I2(n9231), .I3(n11006), .O(n11012) );
  AN2HHD U13716 ( .I1(n11531), .I2(n12480), .O(n10992) );
  OR2KHD U13717 ( .I1(n9232), .I2(n9563), .O(n13408) );
  ND2HHD U13718 ( .I1(n11142), .I2(n9237), .O(n11279) );
  ND2HHD U13719 ( .I1(n9072), .I2(n11439), .O(n11301) );
  ND2KHD U13720 ( .I1(n9626), .I2(n11176), .O(n9237) );
  ND3CHD U13721 ( .I1(n11185), .I2(n11184), .I3(n9238), .O(n11186) );
  ND3EHD U13722 ( .I1(n9679), .I2(n13439), .I3(n9239), .O(n12965) );
  ND3EHD U13723 ( .I1(n8395), .I2(n9241), .I3(n13672), .O(n13676) );
  OAI12CHD U13724 ( .B1(n9243), .B2(n13039), .A1(n13426), .O(n9242) );
  ND2HHD U13725 ( .I1(n13031), .I2(n9252), .O(n9251) );
  OR3HHD U13726 ( .I1(n9232), .I2(n13020), .I3(n9672), .O(n13467) );
  XOR2EHD U13727 ( .I1(n13741), .I2(n9255), .O(n13730) );
  NR2IHD U13728 ( .I1(n8179), .I2(n9256), .O(n10567) );
  ND2HHD U13729 ( .I1(n9531), .I2(n11438), .O(n10569) );
  ND2HHD U13730 ( .I1(n11440), .I2(n9531), .O(n12493) );
  ND3EHD U13731 ( .I1(n12512), .I2(n9260), .I3(n9258), .O(n12515) );
  ND2HHD U13732 ( .I1(n9594), .I2(n9262), .O(n10278) );
  AN3HHD U13733 ( .I1(n8256), .I2(n12490), .I3(n9263), .O(n9262) );
  NR2CHD U13734 ( .I1(n9223), .I2(n12488), .O(n9263) );
  ND2KHD U13735 ( .I1(n9087), .I2(n9800), .O(n12500) );
  OR2B1CHD U13736 ( .I1(n6567), .B1(n10712), .O(n10713) );
  ND2HHD U13737 ( .I1(n9087), .I2(n6873), .O(n11529) );
  ND2KHD U13738 ( .I1(n9266), .I2(n9264), .O(n10208) );
  ND2HHD U13739 ( .I1(n9271), .I2(n9265), .O(n9264) );
  ND2HHD U13740 ( .I1(n9660), .I2(n9987), .O(n9271) );
  XNR2KHD U13741 ( .I1(n9923), .I2(n7868), .O(n14367) );
  ND2HHD U13742 ( .I1(n10559), .I2(_i_CLEFIA128_state_reg _1), .O(n9277) );
  NR2IHD U13743 ( .I1(n10557), .I2(n14707), .O(n9278) );
  AN2HHD U13744 ( .I1(n9285), .I2(n9279), .O(n9557) );
  OAI12CHD U13745 ( .B1(n12961), .B2(n9280), .A1(n13431), .O(n9279) );
  INVCKGHD U13746 ( .I(n9387), .O(n9283) );
  OAI13BHD U13747 ( .B1(n12434), .B2(n13436), .B3(n9286), .A1(n8264), .O(n9285) );
  NR2IHD U13748 ( .I1(n12420), .I2(n12421), .O(n13014) );
  ND3EHD U13749 ( .I1(n8402), .I2(n8234), .I3(n12433), .O(n13436) );
  ND3EHD U13750 ( .I1(n9293), .I2(n9290), .I3(n8239), .O(n9289) );
  NR2GHD U13751 ( .I1(n9291), .I2(n11305), .O(n9290) );
  ND2HHD U13752 ( .I1(n11306), .I2(n11307), .O(n11000) );
  ND2KHD U13753 ( .I1(n8209), .I2(n7810), .O(n9300) );
  XOR2HHD U13754 ( .I1(n8309), .I2(n13717), .O(n9914) );
  ND2HHD U13755 ( .I1(n9303), .I2(n9306), .O(n13717) );
  NR2GHD U13756 ( .I1(n9304), .I2(n9305), .O(n9303) );
  OA13EHD U13757 ( .B1(n12647), .B2(n12649), .B3(n12648), .A1(n12646), .O(n9304) );
  NR2GHD U13758 ( .I1(n9308), .I2(n9307), .O(n9306) );
  ND2HHD U13759 ( .I1(n13829), .I2(n9309), .O(n13525) );
  ND2HHD U13760 ( .I1(n13539), .I2(n8325), .O(n13540) );
  ND2HHD U13761 ( .I1(n8916), .I2(n7420), .O(n9310) );
  AN2HHD U13762 ( .I1(n12338), .I2(n13420), .O(n9311) );
  ND2HHD U13763 ( .I1(n12181), .I2(n13471), .O(n9314) );
  ND3EHD U13764 ( .I1(n9319), .I2(n9323), .I3(n9318), .O(n9317) );
  INVDHD U13765 ( .I(n9324), .O(n9319) );
  ND2HHD U13766 ( .I1(n9324), .I2(n11986), .O(n9322) );
  ND3EHD U13767 ( .I1(n8403), .I2(n12715), .I3(n9459), .O(n9325) );
  ND2KHD U13768 ( .I1(n11713), .I2(n7386), .O(n11814) );
  ND2HHD U13769 ( .I1(n9328), .I2(n8354), .O(n6184) );
  AN2HHD U13770 ( .I1(n13428), .I2(n13424), .O(n9338) );
  NR2CHD U13771 ( .I1(n13375), .I2(n13374), .O(n13428) );
  NR2EHD U13772 ( .I1(n12175), .I2(n9340), .O(n12176) );
  ND2CHD U13773 ( .I1(n8412), .I2(n9339), .O(n13551) );
  ND2HHD U13774 ( .I1(n9341), .I2(n9632), .O(n12442) );
  NR2GHD U13775 ( .I1(n11931), .I2(n11932), .O(n9343) );
  ND2KHD U13776 ( .I1(n7161), .I2(n10179), .O(n9344) );
  ND3EHD U13777 ( .I1(n11229), .I2(n11220), .I3(n9344), .O(n11203) );
  ND3EHD U13778 ( .I1(n12811), .I2(n12806), .I3(n8323), .O(n9346) );
  NR2IHD U13779 ( .I1(n9352), .I2(n9353), .O(n12725) );
  XOR2HHD U13780 ( .I1(DOUT_71), .I2(n9370), .O(n9362) );
  ND3EHD U13781 ( .I1(n13492), .I2(n13493), .I3(n9363), .O(n10193) );
  NR2IHD U13782 ( .I1(n8212), .I2(n10363), .O(n9366) );
  ND2KHD U13783 ( .I1(n11766), .I2(n7907), .O(n9742) );
  ND2KHD U13784 ( .I1(n9368), .I2(n9369), .O(n9370) );
  AN2HHD U13785 ( .I1(n9372), .I2(n13499), .O(n9368) );
  OAI12CHD U13786 ( .B1(n13475), .B2(n13476), .A1(n14049), .O(n9372) );
  XNR2KHD U13787 ( .I1(n8405), .I2(n9376), .O(n12846) );
  ND3EHD U13788 ( .I1(n10405), .I2(n10406), .I3(_i_CLEFIA128_state_reg _1), .O(n9376) );
  AO12EHD U13789 ( .B1(n12841), .B2(n9377), .A1(n12840), .O(n12885) );
  BUFQHD U13790 ( .I(n10427), .O(n9383) );
  ND2DHD U13791 ( .I1(n9389), .I2(n8293), .O(n9440) );
  INVLHD U13792 ( .I(_i_CLEFIA128_keyL _116), .O(n14499) );
  ND2KHD U13793 ( .I1(n8039), .I2(_i_CLEFIA128_keyK _52), .O(n9391) );
  ND3EHD U13794 ( .I1(n9395), .I2(n9394), .I3(n9393), .O(n9392) );
  ND2HHD U13795 ( .I1(n14377), .I2(_i_CLEFIA128_keyL _116), .O(n9396) );
  ND2KHD U13796 ( .I1(n8214), .I2(n12226), .O(n9398) );
  NR2GHD U13797 ( .I1(n9401), .I2(n9399), .O(n14090) );
  OA13EHD U13798 ( .B1(n9402), .B2(n9445), .B3(n14050), .A1(n14049), .O(n9401));
  ND2HHD U13799 ( .I1(n8238), .I2(n8332), .O(n9402) );
  MUX2HHD U13800 ( .A(n14093), .B(n14092), .S(n14613), .O(n14101) );
  XOR2HHD U13801 ( .I1(n14091), .I2(n9407), .O(n14613) );
  ND2KHD U13802 ( .I1(n10473), .I2(n7675), .O(n11511) );
  ND2KHD U13803 ( .I1(n12610), .I2(n9423), .O(n12658) );
  NR2GHD U13804 ( .I1(n9427), .I2(n9426), .O(n9425) );
  ND2HHD U13805 ( .I1(n11236), .I2(n11070), .O(n9427) );
  ND2HHD U13806 ( .I1(n9609), .I2(n6930), .O(n9429) );
  ND2HHD U13807 ( .I1(n8196), .I2(n9435), .O(n11787) );
  NR2IHD U13808 ( .I1(n12214), .I2(n11908), .O(n9436) );
  ND2HHD U13809 ( .I1(n8232), .I2(n12847), .O(n9441) );
  XOR2HHD U13810 ( .I1(n9797), .I2(n9657), .O(n13753) );
  ND3CHD U13811 ( .I1(n11164), .I2(n11178), .I3(n6520), .O(n11165) );
  ND2KHD U13812 ( .I1(n12424), .I2(n9449), .O(n13024) );
  ND2KHD U13813 ( .I1(n9676), .I2(n9449), .O(n13459) );
  ND2KHD U13814 ( .I1(n8214), .I2(n9449), .O(n12419) );
  ND2KHD U13815 ( .I1(n13442), .I2(n9449), .O(n10295) );
  NR2IHD U13816 ( .I1(n10106), .I2(n9458), .O(n12411) );
  INVCKGHD U13817 ( .I(n10034), .O(n9459) );
  OAI22CHD U13818 ( .A1(n7128), .A2(n9613), .B1(n10804), .B2(n10803), .O(n10805) );
  ND3EHD U13819 ( .I1(n11133), .I2(n9461), .I3(n11188), .O(n11134) );
  AN2HHD U13820 ( .I1(n11522), .I2(n12486), .O(n9461) );
  OAI112BHD U13821 ( .C1(n15178), .C2(n8389), .A1(n9464), .B1(n14003), .O(n6136) );
  ND2HHD U13822 ( .I1(n15178), .I2(n8270), .O(n9464) );
  XNR2KHD U13823 ( .I1(n14006), .I2(n9465), .O(n15178) );
  XNR2HHD U13824 ( .I1(n13501), .I2(n13500), .O(n9465) );
  ND2HHD U13825 ( .I1(n10893), .I2(n6734), .O(n9467) );
  XNR2KHD U13826 ( .I1(n10503), .I2(n9469), .O(n12768) );
  NR2CHD U13827 ( .I1(n9270), .I2(n9471), .O(n9470) );
  XOR2HHD U13828 ( .I1(n12014), .I2(n9475), .O(n12054) );
  ND2HHD U13829 ( .I1(n8375), .I2(n9476), .O(n9475) );
  ND2KHD U13830 ( .I1(n12173), .I2(n9479), .O(n9741) );
  ND2HHD U13831 ( .I1(n11818), .I2(n9183), .O(n13088) );
  OR3HHD U13832 ( .I1(n9487), .I2(n9486), .I3(n9485), .O(n9483) );
  NR2GHD U13833 ( .I1(n9491), .I2(n13097), .O(n9490) );
  AN2HHD U13834 ( .I1(n14080), .I2(n12208), .O(n9492) );
  ND2KHD U13835 ( .I1(_i_CLEFIA128_keyK _61), .I2(n8797), .O(n9494) );
  XOR2HHD U13836 ( .I1(n8762), .I2(n9495), .O(n10042) );
  ND3EHD U13837 ( .I1(n13477), .I2(n9508), .I3(n9512), .O(n9650) );
  NR2GHD U13838 ( .I1(n9503), .I2(n9504), .O(n13477) );
  ND2HHD U13839 ( .I1(n8362), .I2(n8253), .O(n9503) );
  ND3EHD U13840 ( .I1(n9506), .I2(n8383), .I3(n9505), .O(n9504) );
  ND2HHD U13841 ( .I1(n9511), .I2(n9510), .O(n9509) );
  NR2CHD U13842 ( .I1(n9513), .I2(n9367), .O(n9512) );
  OR3HHD U13843 ( .I1(n9515), .I2(n9514), .I3(n13252), .O(n9513) );
  ND3EHD U13844 ( .I1(n14071), .I2(n14043), .I3(n9185), .O(n9515) );
  ND3EHD U13845 ( .I1(n11633), .I2(n9517), .I3(n11632), .O(n11637) );
  ND3EHD U13846 ( .I1(n9517), .I2(n11850), .I3(n11851), .O(n11853) );
  ND2CHD U13847 ( .I1(n9604), .I2(n7810), .O(n13841) );
  ND2KHD U13848 ( .I1(n9811), .I2(n7810), .O(n13541) );
  OR3CHD U13849 ( .I1(n13679), .I2(n13678), .I3(n9525), .O(n13687) );
  NR2GHD U13850 ( .I1(_i_CLEFIA128_keyK _73), .I2(n9528), .O(n9527) );
  INVGHD U13851 ( .I(n9530), .O(n10084) );
  BUFQHD U13852 ( .I(n10567), .O(n11274) );
  ND2DHD U13853 ( .I1(n11816), .I2(n13821), .O(n11817) );
  INVGHD U13854 ( .I(n10130), .O(n12044) );
  ND3EHD U13855 ( .I1(n12631), .I2(n12630), .I3(n12629), .O(n12632) );
  INVGHD U13856 ( .I(n11203), .O(n9533) );
  AN2HHD U13857 ( .I1(n11315), .I2(n11314), .O(n11316) );
  AN2HHD U13858 ( .I1(n13366), .I2(n12431), .O(n11949) );
  BUFQHD U13859 ( .I(n11334), .O(n9898) );
  BUFQHD U13860 ( .I(n11895), .O(n11948) );
  ND2HHD U13861 ( .I1(_i_CLEFIA128_keyK _60), .I2(_i_CLEFIA128_keyL _60), .O(n11585) );
  ND2HHD U13862 ( .I1(n10978), .I2(n11531), .O(n11157) );
  ND2HHD U13863 ( .I1(n9804), .I2(n9805), .O(n14327) );
  ND2HHD U13864 ( .I1(n11287), .I2(n11290), .O(n10724) );
  ND2HHD U13865 ( .I1(n11015), .I2(n11349), .O(n9795) );
  MUX2HHD U13866 ( .A(n13940), .B(n13939), .S(n15377), .O(n13948) );
  ND2HHD U13867 ( .I1(n12610), .I2(n11254), .O(n11065) );
  XOR2HHD U13868 ( .I1(DOUT_31), .I2(n9960), .O(n9544) );
  ND2HHD U13869 ( .I1(n12792), .I2(n10207), .O(n12851) );
  INVKHD U13870 ( .I(n9755), .O(n14621) );
  ND2HHD U13871 ( .I1(n13440), .I2(n13400), .O(n12440) );
  ND2KHD U13872 ( .I1(n8214), .I2(n12327), .O(n13440) );
  NR2GHD U13873 ( .I1(n13583), .I2(n13584), .O(n13626) );
  ND3EHD U13874 ( .I1(n11949), .I2(n9574), .I3(n13019), .O(n11951) );
  OAI112BHD U13875 ( .C1(n15435), .C2(n13769), .A1(n9545), .B1(n13776), .O(n6135) );
  ND2HHD U13876 ( .I1(n15435), .I2(n8271), .O(n9545) );
  ND3EHD U13877 ( .I1(n9546), .I2(n9999), .I3(n8300), .O(n6201) );
  ND2HHD U13878 ( .I1(n12743), .I2(n12586), .O(n11383) );
  INVNHD U13879 ( .I(n12914), .O(n10131) );
  ND3EHD U13880 ( .I1(n9552), .I2(n13250), .I3(n13249), .O(n9551) );
  ND2HHD U13881 ( .I1(n9766), .I2(n10632), .O(n11234) );
  BUFQHD U13882 ( .I(n10424), .O(n12829) );
  ND2HHD U13883 ( .I1(n11902), .I2(n11901), .O(n13381) );
  AN3HHD U13884 ( .I1(n12620), .I2(n8235), .I3(n11221), .O(n12603) );
  AN2HHD U13885 ( .I1(n12621), .I2(n12537), .O(n11255) );
  BUFEHD U13886 ( .I(n8199), .O(n9561) );
  AN2HHD U13887 ( .I1(n11230), .I2(n11216), .O(n12605) );
  ND3EHD U13888 ( .I1(n13477), .I2(n13240), .I3(n13239), .O(n13242) );
  INVNHD U13889 ( .I(n9562), .O(n9766) );
  ND3CHD U13890 ( .I1(n11740), .I2(n8253), .I3(n13222), .O(n11741) );
  ND2HHD U13891 ( .I1(n6753), .I2(n13440), .O(n9563) );
  NR2EHD U13892 ( .I1(n12146), .I2(n12147), .O(n12148) );
  ND2HHD U13893 ( .I1(n9684), .I2(n10969), .O(n12866) );
  ND2HHD U13894 ( .I1(n12436), .I2(n9847), .O(n13388) );
  ND2KHD U13895 ( .I1(n10225), .I2(n11612), .O(n11839) );
  INVGHD U13896 ( .I(n10450), .O(n9590) );
  NR2GHD U13897 ( .I1(n13435), .I2(n12990), .O(n12992) );
  XOR2HHD U13898 ( .I1(n10042), .I2(n14331), .O(n9571) );
  INVGHD U13899 ( .I(n13253), .O(n11750) );
  XNR2KHD U13900 ( .I1(n14194), .I2(n9571), .O(n14601) );
  XNR3EHD U13901 ( .I1(n14015), .I2(n13741), .I3(n14489), .O(n14144) );
  ND3EHD U13902 ( .I1(n11972), .I2(n11971), .I3(n11970), .O(n9572) );
  ND2HHD U13903 ( .I1(n11232), .I2(n11201), .O(n10234) );
  BUFKHD U13904 ( .I(n10295), .O(n9574) );
  ND2HHD U13905 ( .I1(n12538), .I2(n10776), .O(n10646) );
  ND2HHD U13906 ( .I1(n13072), .I2(n14078), .O(n13073) );
  INVGHD U13907 ( .I(n9770), .O(n12046) );
  ND2KHD U13908 ( .I1(n12900), .I2(n12383), .O(n13191) );
  ND2HHD U13909 ( .I1(n9586), .I2(_i_CLEFIA128_keyL _44), .O(n9660) );
  AN2HHD U13910 ( .I1(n13577), .I2(n13125), .O(n12048) );
  ND2HHD U13911 ( .I1(n12749), .I2(n11323), .O(n11474) );
  NR2IHD U13912 ( .I1(n9969), .I2(n11156), .O(n11306) );
  ND2KHD U13913 ( .I1(n12327), .I2(n11948), .O(n12364) );
  ND2HHD U13914 ( .I1(n12968), .I2(n12970), .O(n12348) );
  OA112EHD U13915 ( .C1(n13219), .C2(n13218), .A1(n13217), .B1(n6632), .O(n13221) );
  INVCKIHD U13916 ( .I(n12305), .O(n11774) );
  ND2KHD U13917 ( .I1(n11906), .I2(n7032), .O(n12988) );
  BUFEHD U13918 ( .I(n12477), .O(n9594) );
  ND3EHD U13919 ( .I1(n11344), .I2(n12777), .I3(n11343), .O(n11345) );
  ND2HHD U13920 ( .I1(n9895), .I2(n8284), .O(n9719) );
  ND2HHD U13921 ( .I1(n10798), .I2(n9709), .O(n11242) );
  OR2KHD U13922 ( .I1(n12334), .I2(n9672), .O(n9990) );
  OR3HHD U13923 ( .I1(n12918), .I2(n12396), .I3(n13173), .O(n12397) );
  OR3HHD U13924 ( .I1(n10782), .I2(n10863), .I3(n10781), .O(n10788) );
  ND2HHD U13925 ( .I1(n12521), .I2(n12522), .O(n11058) );
  ND2HHD U13926 ( .I1(n13908), .I2(n13907), .O(n6109) );
  ND2HHD U13927 ( .I1(n8278), .I2(n11489), .O(n9600) );
  XNR2HHD U13928 ( .I1(n13896), .I2(n13895), .O(n13898) );
  AN2HHD U13929 ( .I1(n13478), .I2(n13085), .O(n14046) );
  ND3EHD U13930 ( .I1(n9623), .I2(n12443), .I3(n9722), .O(n12444) );
  BUFQHD U13931 ( .I(n10570), .O(n10599) );
  AN3HHD U13932 ( .I1(n9873), .I2(n13447), .I3(n12419), .O(n13031) );
  OR3HHD U13933 ( .I1(n11936), .I2(n12238), .I3(n12967), .O(n12322) );
  OR3HHD U13934 ( .I1(n11224), .I2(n10836), .I3(n10835), .O(n10838) );
  AN2HHD U13935 ( .I1(n13841), .I2(n9741), .O(n13843) );
  OR3HHD U13936 ( .I1(n10538), .I2(n10536), .I3(n10537), .O(n12761) );
  ND3EHD U13937 ( .I1(n10244), .I2(n10242), .I3(n10464), .O(n10058) );
  AN2HHD U13938 ( .I1(n12419), .I2(n13398), .O(n12369) );
  BUFEHD U13939 ( .I(n11930), .O(n9609) );
  INVJHD U13940 ( .I(n12468), .O(n9969) );
  ND2KHD U13941 ( .I1(n8180), .I2(n9050), .O(n11368) );
  INVGHD U13942 ( .I(n11712), .O(n9845) );
  ND2HHD U13943 ( .I1(n12087), .I2(n12088), .O(n11712) );
  NR2EHD U13944 ( .I1(n12800), .I2(n12691), .O(n12698) );
  AN2HHD U13945 ( .I1(n13398), .I2(n12219), .O(n12220) );
  OR3HHD U13946 ( .I1(n13124), .I2(n13123), .I3(n13605), .O(n10132) );
  ND2HHD U13947 ( .I1(n9611), .I2(n9986), .O(n9985) );
  INVGHD U13948 ( .I(n12571), .O(n12572) );
  ND2KHD U13949 ( .I1(n9597), .I2(n9186), .O(n13102) );
  OR3HHD U13950 ( .I1(n13455), .I2(n13456), .I3(n13454), .O(n13468) );
  ND3EHD U13951 ( .I1(n11456), .I2(n11457), .I3(n12467), .O(n11458) );
  NR2GHD U13952 ( .I1(n11162), .I2(n11163), .O(n11457) );
  NR2CHD U13953 ( .I1(n15513), .I2(n14766), .O(n14007) );
  ND2KHD U13954 ( .I1(n7039), .I2(n9050), .O(n12729) );
  ND2HHD U13955 ( .I1(n13681), .I2(n12080), .O(n13670) );
  INVQHD U13956 ( .I(n9613), .O(n9730) );
  AN2HHD U13957 ( .I1(n12062), .I2(n12063), .O(n13634) );
  XNR2KHD U13958 ( .I1(n13911), .I2(n10229), .O(n13926) );
  NR2IHD U13959 ( .I1(n13617), .I2(n9614), .O(n13179) );
  NR2IHD U13960 ( .I1(n12224), .I2(n13449), .O(n12981) );
  ND2HHD U13961 ( .I1(n11552), .I2(n10588), .O(n10589) );
  BUFKHD U13962 ( .I(n12582), .O(n9682) );
  OA13EHD U13963 ( .B1(n12116), .B2(n12115), .B3(n13636), .A1(n13585), .O(n12137) );
  INVDHD U13964 ( .I(n12057), .O(n9736) );
  ND2HHD U13965 ( .I1(n13474), .I2(n11835), .O(n11836) );
  ND3EHD U13966 ( .I1(n11267), .I2(n11266), .I3(n12615), .O(n11268) );
  ND2HHD U13967 ( .I1(n10783), .I2(n11216), .O(n10870) );
  ND3EHD U13968 ( .I1(n9617), .I2(n13049), .I3(n13048), .O(n6140) );
  AN2HHD U13969 ( .I1(n8408), .I2(n13014), .O(n9623) );
  ND2KHD U13970 ( .I1(n10599), .I2(n12484), .O(n11192) );
  NR2IHD U13971 ( .I1(n11903), .I2(n12975), .O(n9918) );
  OR3HHD U13972 ( .I1(n10585), .I2(n10584), .I3(n11276), .O(n11137) );
  AN2HHD U13973 ( .I1(n12549), .I2(n12550), .O(n9624) );
  ND3EHD U13974 ( .I1(n11513), .I2(n12585), .I3(n12729), .O(n11514) );
  ND2HHD U13975 ( .I1(n8432), .I2(n12278), .O(n13635) );
  ND2HHD U13976 ( .I1(n11213), .I2(n11214), .O(n11215) );
  OR3HHD U13977 ( .I1(n12911), .I2(n12941), .I3(n9629), .O(n12912) );
  BUFKHD U13978 ( .I(n9847), .O(n9846) );
  INVNHD U13979 ( .I(n11548), .O(n9964) );
  ND3EHD U13980 ( .I1(n8245), .I2(n9630), .I3(n6932), .O(n13064) );
  ND2KHD U13981 ( .I1(n11415), .I2(n10089), .O(n13741) );
  ND3EHD U13982 ( .I1(n13119), .I2(n13120), .I3(n13118), .O(n13157) );
  INVGHD U13983 ( .I(n12614), .O(n10016) );
  ND2HHD U13984 ( .I1(n15307), .I2(n11130), .O(n14676) );
  AN2HHD U13985 ( .I1(n13021), .I2(n12427), .O(n13406) );
  ND2HHD U13986 ( .I1(n7703), .I2(n7907), .O(n13077) );
  BUFKHD U13987 ( .I(n10229), .O(n9637) );
  ND3EHD U13988 ( .I1(n11743), .I2(n11742), .I3(n13246), .O(n11749) );
  ND3EHD U13989 ( .I1(n13491), .I2(n13062), .I3(n11747), .O(n12188) );
  AN2HHD U13990 ( .I1(n10797), .I2(n10873), .O(n10799) );
  INVNHD U13991 ( .I(n10074), .O(n12743) );
  ND2HHD U13992 ( .I1(n13582), .I2(n13628), .O(n12052) );
  ND3EHD U13993 ( .I1(n11941), .I2(n9641), .I3(n11940), .O(n11946) );
  AN3HHD U13994 ( .I1(n13366), .I2(n13021), .I3(n13419), .O(n12225) );
  INVGHD U13995 ( .I(n13591), .O(n13115) );
  ND2HHD U13996 ( .I1(n12917), .I2(n13628), .O(n13124) );
  AN2HHD U13997 ( .I1(n12622), .I2(n12521), .O(n10785) );
  ND2KHD U13998 ( .I1(n13442), .I2(n12251), .O(n13419) );
  NR2GHD U13999 ( .I1(n11755), .I2(n8794), .O(n11821) );
  INVGHD U14000 ( .I(n11989), .O(n10112) );
  ND3EHD U14001 ( .I1(n8401), .I2(n13111), .I3(n13110), .O(n10154) );
  ND3EHD U14002 ( .I1(n12755), .I2(n12749), .I3(n8366), .O(n12756) );
  ND2HHD U14003 ( .I1(n13396), .I2(n12364), .O(n13446) );
  OR2EHD U14004 ( .I1(n13496), .I2(n13495), .O(n13497) );
  ND3EHD U14005 ( .I1(n8202), .I2(n11233), .I3(n11234), .O(n11060) );
  ND2KHD U14006 ( .I1(n6872), .I2(n7809), .O(n13837) );
  NR2EHD U14007 ( .I1(n12334), .I2(n12965), .O(n13404) );
  INVGHD U14008 ( .I(n12319), .O(n9814) );
  ND3EHD U14009 ( .I1(n9652), .I2(n11003), .I3(n11002), .O(n10184) );
  NR2IHD U14010 ( .I1(n13639), .I2(n13638), .O(n13640) );
  OR3HHD U14011 ( .I1(n12503), .I2(n11462), .I3(n11461), .O(n11468) );
  ND3EHD U14012 ( .I1(n10245), .I2(n10462), .I3(_i_CLEFIA128_state_reg _1), .O(n9654) );
  ND3EHD U14013 ( .I1(n11761), .I2(n13076), .I3(n13084), .O(n13238) );
  ND3EHD U14014 ( .I1(n6707), .I2(n13220), .I3(n13221), .O(n13227) );
  ND2HHD U14015 ( .I1(n15307), .I2(n15500), .O(n14673) );
  ND2HHD U14016 ( .I1(_i_CLEFIA128_keyK _50), .I2(_i_CLEFIA128_keyL _50), .O(n11671) );
  NR2GHD U14017 ( .I1(n13235), .I2(n11657), .O(n11743) );
  ND2HHD U14018 ( .I1(n13573), .I2(n12287), .O(n12289) );
  XOR2HHD U14019 ( .I1(_i_CLEFIA128_keyL _124), .I2(n11586), .O(n11588) );
  ND2HHD U14020 ( .I1(n10760), .I2(n8938), .O(n10893) );
  OR3HHD U14021 ( .I1(n12381), .I2(n12380), .I3(n12379), .O(n12382) );
  ND2HHD U14022 ( .I1(n7041), .I2(n9811), .O(n12153) );
  ND2HHD U14023 ( .I1(n9991), .I2(n10436), .O(n10437) );
  ND2KHD U14024 ( .I1(n8320), .I2(n12439), .O(n13435) );
  ND3EHD U14025 ( .I1(n10880), .I2(n10878), .I3(n10879), .O(n9665) );
  BUFKHD U14026 ( .I(n12769), .O(n9666) );
  ND2HHD U14027 ( .I1(n11069), .I2(n12521), .O(n10795) );
  AN2HHD U14028 ( .I1(n12730), .I2(n12729), .O(n12732) );
  ND2KHD U14029 ( .I1(n9699), .I2(n8185), .O(n9886) );
  ND2KHD U14030 ( .I1(n9699), .I2(n12383), .O(n10080) );
  OAI112BHD U14031 ( .C1(n14575), .C2(n14157), .A1(n9670), .B1(n14164), .O(n6141) );
  ND2HHD U14032 ( .I1(n14575), .I2(n8272), .O(n9670) );
  XOR2HHD U14033 ( .I1(n9705), .I2(n9776), .O(n14768) );
  OA13EHD U14034 ( .B1(n11115), .B2(n11357), .B3(n11116), .A1(n11479), .O(n11127) );
  ND2HHD U14035 ( .I1(n12988), .I2(n13396), .O(n12233) );
  ND2KHD U14036 ( .I1(n9964), .I2(n7671), .O(n12454) );
  ND2KHD U14037 ( .I1(n9597), .I2(n7907), .O(n14056) );
  ND2HHD U14038 ( .I1(n12730), .I2(n11512), .O(n12744) );
  ND2KHD U14039 ( .I1(n9694), .I2(n9049), .O(n11340) );
  ND2KHD U14040 ( .I1(n6873), .I2(n12498), .O(n11155) );
  ND2HHD U14041 ( .I1(n13200), .I2(n7031), .O(n13201) );
  BUFEHD U14042 ( .I(n9456), .O(n9674) );
  ND3EHD U14043 ( .I1(n9862), .I2(n9865), .I3(n12997), .O(n10159) );
  ND2KHD U14044 ( .I1(n12125), .I2(n8185), .O(n12905) );
  ND2HHD U14045 ( .I1(_i_CLEFIA128_keyK _25), .I2(_i_CLEFIA128_keyL _25), .O(n10322) );
  ND2HHD U14046 ( .I1(_i_CLEFIA128_keyK _13), .I2(_i_CLEFIA128_keyL _13), .O(n10414) );
  ND2HHD U14047 ( .I1(n13764), .I2(n13763), .O(n6118) );
  AN2HHD U14048 ( .I1(n12410), .I2(n12436), .O(n13441) );
  AN3B1HHD U14049 ( .I1(n13031), .I2(n13386), .B1(n13029), .O(n13370) );
  XNR2KHD U14050 ( .I1(n9816), .I2(n14215), .O(n14171) );
  ND3EHD U14051 ( .I1(n13448), .I2(n11937), .I3(n9026), .O(n11938) );
  OR2KHD U14052 ( .I1(n11129), .I2(n15449), .O(n15448) );
  OR3HHD U14053 ( .I1(n12994), .I2(n12993), .I3(n13039), .O(n12995) );
  INVMHD U14054 ( .I(_i_CLEFIA128_keyK _69), .O(n14242) );
  ND3EHD U14055 ( .I1(n13024), .I2(n13000), .I3(n12963), .O(n13017) );
  INVCKGHD U14056 ( .I(n13050), .O(n12996) );
  BUFQHD U14057 ( .I(n12056), .O(n12291) );
  INVGHD U14058 ( .I(n7128), .O(n10271) );
  AN2HHD U14059 ( .I1(n10905), .I2(n12868), .O(n10810) );
  ND2KHD U14060 ( .I1(n11818), .I2(n8210), .O(n14080) );
  OR3HHD U14061 ( .I1(n10936), .I2(n10742), .I3(n12665), .O(n10743) );
  ND2KHD U14062 ( .I1(n10123), .I2(n9684), .O(n12867) );
  ND2KHD U14063 ( .I1(n12876), .I2(n8193), .O(n10967) );
  ND3EHD U14064 ( .I1(n11770), .I2(n11769), .I3(n11768), .O(n11771) );
  ND2KHD U14065 ( .I1(n8183), .I2(n12915), .O(n13130) );
  AN2KHD U14066 ( .I1(n13241), .I2(n13233), .O(n14049) );
  OA22HHD U14067 ( .A1(n10654), .A2(n10655), .B1(n10656), .B2(n10683), .O(n10687) );
  MUX2HHD U14068 ( .A(n13872), .B(n13871), .S(n15269), .O(n13880) );
  ND2KHD U14069 ( .I1(n11648), .I2(n7044), .O(n11593) );
  ND2KHD U14070 ( .I1(n11284), .I2(n11438), .O(n11159) );
  ND3EHD U14071 ( .I1(n8246), .I2(n9688), .I3(n8436), .O(n9968) );
  AN2HHD U14072 ( .I1(n10644), .I2(n10384), .O(n9690) );
  ND2KHD U14073 ( .I1(n9559), .I2(n9383), .O(n9916) );
  ND3EHD U14074 ( .I1(n10204), .I2(n8311), .I3(n10203), .O(n6168) );
  ND3EHD U14075 ( .I1(n11656), .I2(n11655), .I3(n14065), .O(n9692) );
  ND2KHD U14076 ( .I1(n10179), .I2(n10011), .O(n9709) );
  INVCKGHD U14077 ( .I(n12668), .O(n10764) );
  OR3HHD U14078 ( .I1(n11620), .I2(n11619), .I3(n11618), .O(n11624) );
  NR2EHD U14079 ( .I1(n12388), .I2(n12262), .O(n12263) );
  ND3EHD U14080 ( .I1(n8798), .I2(n14419), .I3(_i_CLEFIA128_rndcnt_reg _4), .O(n13287) );
  ND3EHD U14081 ( .I1(n12200), .I2(n12199), .I3(n11831), .O(n9696) );
  OAI112BHD U14082 ( .C1(n15193), .C2(n14117), .A1(n9698), .B1(n14124), .O(n6150) );
  AN3HHD U14083 ( .I1(n13372), .I2(n12427), .I3(n9847), .O(n12970) );
  ND2KHD U14084 ( .I1(n10059), .I2(n10058), .O(n10481) );
  ND3EHD U14085 ( .I1(n9982), .I2(n9984), .I3(n9983), .O(n9701) );
  ND2KHD U14086 ( .I1(n7398), .I2(n12561), .O(n11503) );
  BUFKHD U14087 ( .I(n7955), .O(n9705) );
  ND2KHD U14088 ( .I1(n12190), .I2(n8204), .O(n14082) );
  XNR3EHD U14089 ( .I1(n9710), .I2(n14005), .I3(n14006), .O(n9778) );
  ND3EHD U14090 ( .I1(n10673), .I2(n9648), .I3(n11250), .O(n10362) );
  ND2KHD U14091 ( .I1(n12517), .I2(n10011), .O(n11221) );
  ND2HHD U14092 ( .I1(n11269), .I2(n11268), .O(n11270) );
  ND3EHD U14093 ( .I1(n12602), .I2(n12650), .I3(n12601), .O(n12608) );
  NR2IHD U14094 ( .I1(n8212), .I2(n10332), .O(n10324) );
  ND3EHD U14095 ( .I1(n11308), .I2(n11307), .I3(n11306), .O(n11536) );
  OR3HHD U14096 ( .I1(n12222), .I2(n12223), .I3(n12221), .O(n10100) );
  ND3EHD U14097 ( .I1(n13400), .I2(n12988), .I3(n13459), .O(n12223) );
  AN3HHD U14098 ( .I1(n11287), .I2(n11288), .I3(n11289), .O(n11291) );
  ND2KHD U14099 ( .I1(n9738), .I2(n9050), .O(n12742) );
  ND3EHD U14100 ( .I1(n10350), .I2(n10351), .I3(_i_CLEFIA128_state_reg _1), .O(n10352) );
  NR2GHD U14101 ( .I1(n11341), .I2(n11392), .O(n11342) );
  OAI112BHD U14102 ( .C1(n15095), .C2(n14203), .A1(n9714), .B1(n14210), .O(n6145) );
  OAI112BHD U14103 ( .C1(n9817), .C2(n14297), .A1(n9715), .B1(n14305), .O(n6137) );
  OAI12CHD U14104 ( .B1(n11125), .B2(n10541), .A1(n12575), .O(n9716) );
  OR3HHD U14105 ( .I1(n11005), .I2(n11004), .I3(n12457), .O(n11006) );
  ND2KHD U14106 ( .I1(n8180), .I2(n9898), .O(n12765) );
  ND3EHD U14107 ( .I1(n13400), .I2(n13366), .I3(n13000), .O(n12345) );
  OAI112BHD U14108 ( .C1(n9895), .C2(n14368), .A1(n9719), .B1(n14375), .O(n6139) );
  XNR2KHD U14109 ( .I1(n13215), .I2(n9978), .O(n14344) );
  ND2KHD U14110 ( .I1(n7038), .I2(n12251), .O(n13396) );
  ND2KHD U14111 ( .I1(n7777), .I2(n10145), .O(n11793) );
  ND2KHD U14112 ( .I1(n11049), .I2(n9898), .O(n12578) );
  NR2GHD U14113 ( .I1(n11666), .I2(n14707), .O(n9721) );
  NR2EHD U14114 ( .I1(n12720), .I2(n10527), .O(n10532) );
  AN2HHD U14115 ( .I1(n12578), .I2(n12577), .O(n12767) );
  ND2HHD U14116 ( .I1(n12743), .I2(n11368), .O(n11351) );
  AN2HHD U14117 ( .I1(n12581), .I2(n11360), .O(n10250) );
  ND2KHD U14118 ( .I1(n8904), .I2(n8180), .O(n11360) );
  AN2HHD U14119 ( .I1(n10043), .I2(n11472), .O(n9725) );
  OR3HHD U14120 ( .I1(n11017), .I2(n11401), .I3(n11016), .O(n11116) );
  ND2HHD U14121 ( .I1(n12558), .I2(n10073), .O(n12568) );
  ND2KHD U14122 ( .I1(n7830), .I2(n7038), .O(n13004) );
  OAI112BHD U14123 ( .C1(n15134), .C2(n11129), .A1(n8244), .B1(n9729), .O(n6176) );
  ND2KHD U14124 ( .I1(n11175), .I2(n8179), .O(n9758) );
  ND2KHD U14125 ( .I1(n8214), .I2(n12251), .O(n13399) );
  OAI12CHD U14126 ( .B1(n13139), .B2(n13140), .A1(n13608), .O(n9732) );
  ND3EHD U14127 ( .I1(n13179), .I2(n12924), .I3(n12387), .O(n12392) );
  AN2HHD U14128 ( .I1(n11776), .I2(n12153), .O(n11777) );
  ND2KHD U14129 ( .I1(n8767), .I2(n9903), .O(n12453) );
  OA12HHD U14130 ( .B1(n14601), .B2(n11129), .A1(n12447), .O(n12593) );
  ND2KHD U14131 ( .I1(n7034), .I2(n8210), .O(n13076) );
  ND2HHD U14132 ( .I1(n8607), .I2(n12765), .O(n11476) );
  XNR2KHD U14133 ( .I1(n11601), .I2(n11600), .O(n13241) );
  ND3EHD U14134 ( .I1(n12003), .I2(n9736), .I3(n13175), .O(n13140) );
  OR3HHD U14135 ( .I1(n10516), .I2(n10517), .I3(n12758), .O(n12573) );
  ND2KHD U14136 ( .I1(n8209), .I2(n7035), .O(n13513) );
  ND3EHD U14137 ( .I1(n10730), .I2(n12690), .I3(n12668), .O(n10734) );
  ND2HHD U14138 ( .I1(n11263), .I2(n11255), .O(n12526) );
  INVGHD U14139 ( .I(n11044), .O(n11500) );
  XNR2KHD U14140 ( .I1(n10496), .I2(n10495), .O(n12747) );
  ND2KHD U14141 ( .I1(n8771), .I2(n9480), .O(n13844) );
  INVNHD U14142 ( .I(n9822), .O(n10051) );
  ND3EHD U14143 ( .I1(n10045), .I2(n10050), .I3(n11230), .O(n11271) );
  INVGHD U14144 ( .I(n7036), .O(n11779) );
  ND2KHD U14145 ( .I1(n11049), .I2(n11335), .O(n11019) );
  ND2KHD U14146 ( .I1(n12327), .I2(n11906), .O(n12338) );
  XNR3EHD U14147 ( .I1(n10262), .I2(n14636), .I3(n9743), .O(n15336) );
  ND3EHD U14148 ( .I1(n6921), .I2(n10786), .I3(n10785), .O(n10787) );
  OR3HHD U14149 ( .I1(n13232), .I2(n13080), .I3(n13079), .O(n13081) );
  ND2KHD U14150 ( .I1(n15367), .I2(n15355), .O(n15365) );
  OAI112BHD U14151 ( .C1(n14621), .C2(n14286), .A1(n9745), .B1(n14294), .O(n6131) );
  ND2HHD U14152 ( .I1(n14621), .I2(n8298), .O(n9745) );
  XOR2HHD U14153 ( .I1(DOUT_72), .I2(n14227), .O(n9746) );
  INVNHD U14154 ( .I(n11680), .O(n10145) );
  ND2HHD U14155 ( .I1(n10052), .I2(n11412), .O(n9748) );
  ND2KHD U14156 ( .I1(n7507), .I2(n10011), .O(n11254) );
  ND3EHD U14157 ( .I1(n12516), .I2(n10641), .I3(n9656), .O(n10656) );
  NR2GHD U14158 ( .I1(n10021), .I2(n10801), .O(n10638) );
  ND2HHD U14159 ( .I1(n13421), .I2(n9679), .O(n12982) );
  OAI112BHD U14160 ( .C1(n10008), .C2(n14185), .A1(n9753), .B1(n14192), .O(n6129) );
  ND2HHD U14161 ( .I1(n10008), .I2(n8274), .O(n9753) );
  ND2KHD U14162 ( .I1(n9917), .I2(n11948), .O(n13022) );
  ND3EHD U14163 ( .I1(n13607), .I2(n12050), .I3(n12051), .O(n12055) );
  ND2KHD U14164 ( .I1(n9897), .I2(n11335), .O(n11512) );
  NR2CHD U14165 ( .I1(n11313), .I2(n9931), .O(n11315) );
  ND2HHD U14166 ( .I1(n12766), .I2(n11358), .O(n11494) );
  ND3EHD U14167 ( .I1(n11317), .I2(n11316), .I3(n11457), .O(n11319) );
  XNR3EHD U14168 ( .I1(DOUT_10), .I2(n14167), .I3(n7789), .O(n9756) );
  ND2KHD U14169 ( .I1(n7864), .I2(n10011), .O(n10847) );
  ND2KHD U14170 ( .I1(n8797), .I2(_i_CLEFIA128_keyK _112), .O(n11670) );
  ND2HHD U14171 ( .I1(n14272), .I2(n14273), .O(n6202) );
  NR2GHD U14172 ( .I1(n12441), .I2(n12442), .O(n12443) );
  ND2KHD U14173 ( .I1(n9917), .I2(n11906), .O(n13460) );
  OAI112BHD U14174 ( .C1(n15152), .C2(n14127), .A1(n9760), .B1(n14134), .O(n6095) );
  ND2HHD U14175 ( .I1(n15152), .I2(n8275), .O(n9760) );
  ND2KHD U14176 ( .I1(n13442), .I2(n9430), .O(n12427) );
  ND2KHD U14177 ( .I1(n9964), .I2(n10600), .O(n11295) );
  OR3HHD U14178 ( .I1(n9946), .I2(n12998), .I3(n9863), .O(n9862) );
  XOR2HHD U14179 ( .I1(_i_CLEFIA128_CON_T_x _0), .I2(DOUT_96), .O(n11989) );
  ND3EHD U14180 ( .I1(n11524), .I2(n11523), .I3(n11525), .O(n11528) );
  ND2KHD U14181 ( .I1(n8797), .I2(_i_CLEFIA128_keyK _37), .O(n11974) );
  OR3HHD U14182 ( .I1(n12808), .I2(n10732), .I3(n10731), .O(n10733) );
  ND2KHD U14183 ( .I1(n9186), .I2(n9628), .O(n14053) );
  OAI112BHD U14184 ( .C1(n14601), .C2(n14276), .A1(n9762), .B1(n14283), .O(n6130) );
  ND2HHD U14185 ( .I1(n14601), .I2(n8276), .O(n9762) );
  ND2HHD U14186 ( .I1(n14197), .I2(n14198), .O(n6185) );
  ND2KHD U14187 ( .I1(n8180), .I2(n8188), .O(n11349) );
  ND2HHD U14188 ( .I1(n14268), .I2(n14269), .O(n6170) );
  NR2IHD U14189 ( .I1(n9456), .I2(n12000), .O(n9887) );
  MUX2HHD U14190 ( .A(n13900), .B(n13899), .S(n15131), .O(n13908) );
  OR3HHD U14191 ( .I1(n12875), .I2(n12836), .I3(n10729), .O(n12860) );
  AN2HHD U14192 ( .I1(n13283), .I2(n13282), .O(n14721) );
  ND2KHD U14193 ( .I1(n9628), .I2(n7907), .O(n13222) );
  AN2KHD U14194 ( .I1(n14431), .I2(n14430), .O(n14432) );
  XOR2HHD U14195 ( .I1(n14015), .I2(n13715), .O(n9958) );
  XNR2KHD U14196 ( .I1(n14031), .I2(n14030), .O(n15449) );
  ND2KHD U14197 ( .I1(n8768), .I2(n10600), .O(n12464) );
  AN2HHD U14198 ( .I1(n8304), .I2(n13386), .O(n11913) );
  XNR2KHD U14199 ( .I1(n10087), .I2(n10086), .O(n15440) );
  OAI112BHD U14200 ( .C1(n15440), .C2(n14018), .A1(n9767), .B1(n14025), .O(n6121) );
  ND2HHD U14201 ( .I1(n14398), .I2(n14397), .O(n6147) );
  ND2KHD U14202 ( .I1(n10318), .I2(n7864), .O(n12522) );
  AN2HHD U14203 ( .I1(n13527), .I2(n13526), .O(n13528) );
  ND3EHD U14204 ( .I1(n13528), .I2(n13529), .I3(n6684), .O(n13534) );
  ND2KHD U14205 ( .I1(n8797), .I2(_i_CLEFIA128_keyK _59), .O(n11581) );
  XOR2HHD U14206 ( .I1(n10147), .I2(n10004), .O(n10003) );
  XOR3EHD U14207 ( .I1(n14170), .I2(DOUT_21), .I3(n14805), .O(n10211) );
  ND3EHD U14208 ( .I1(n13179), .I2(n13148), .I3(n13147), .O(n13149) );
  ND2KHD U14209 ( .I1(n8797), .I2(_i_CLEFIA128_keyK _16), .O(n10114) );
  BUFEHD U14210 ( .I(n6838), .O(n9776) );
  ND2KHD U14211 ( .I1(n12251), .I2(n9676), .O(n12410) );
  ND2KHD U14212 ( .I1(n13442), .I2(n12327), .O(n12431) );
  OA12HHD U14213 ( .B1(n11125), .B2(n11124), .A1(n11500), .O(n11126) );
  ND2HHD U14214 ( .I1(n15481), .I2(n15470), .O(n15479) );
  ND2HHD U14215 ( .I1(n8797), .I2(_i_CLEFIA128_keyK _33), .O(n11977) );
  INVNHD U14216 ( .I(n10191), .O(n11818) );
  ND2HHD U14217 ( .I1(n9780), .I2(n9781), .O(n6217) );
  OA12HHD U14218 ( .B1(n14621), .B2(n15513), .A1(n14200), .O(n9780) );
  ND2HHD U14219 ( .I1(n9779), .I2(n11130), .O(n9781) );
  XOR2HHD U14220 ( .I1(n9839), .I2(n9838), .O(n9836) );
  ND3EHD U14221 ( .I1(n11320), .I2(n11319), .I3(n11318), .O(n9783) );
  ND2HHD U14222 ( .I1(n10467), .I2(_i_CLEFIA128_state_reg _1), .O(n9786) );
  ND2HHD U14223 ( .I1(n12593), .I2(n9788), .O(n6186) );
  ND3EHD U14224 ( .I1(n9793), .I2(n9792), .I3(n9791), .O(n9790) );
  ND2HHD U14225 ( .I1(n14242), .I2(_i_CLEFIA128_keyL _69), .O(n9794) );
  OR3HHD U14226 ( .I1(n11431), .I2(n11448), .I3(n12503), .O(n9899) );
  OR2KHD U14227 ( .I1(n12137), .I2(n9877), .O(n13556) );
  OR2B1CHD U14228 ( .I1(n11685), .B1(n9549), .O(n11683) );
  INVDHD U14229 ( .I(n13805), .O(n9835) );
  ND2HHD U14230 ( .I1(n9837), .I2(n15250), .O(n6321) );
  ND2HHD U14231 ( .I1(n9779), .I2(n7043), .O(n9837) );
  XOR2HHD U14232 ( .I1(n9938), .I2(n14143), .O(n9838) );
  XOR2HHD U14233 ( .I1(n14142), .I2(n14144), .O(n9839) );
  OR3HHD U14234 ( .I1(n11161), .I2(n11160), .I3(n11159), .O(n11162) );
  ND2KHD U14235 ( .I1(n9676), .I2(n12226), .O(n9847) );
  ND3EHD U14236 ( .I1(n13367), .I2(n12976), .I3(n9846), .O(n12977) );
  ND3EHD U14237 ( .I1(n12956), .I2(n12955), .I3(n9846), .O(n12957) );
  ND3EHD U14238 ( .I1(n9850), .I2(n9853), .I3(n12856), .O(n9849) );
  ND3EHD U14239 ( .I1(n9852), .I2(n10824), .I3(n9851), .O(n9850) );
  ND3EHD U14240 ( .I1(n10832), .I2(n10831), .I3(n9854), .O(n9853) );
  OAI12CHD U14241 ( .B1(n9089), .B2(n11129), .A1(n9856), .O(n6189) );
  ND2HHD U14242 ( .I1(n9864), .I2(n13050), .O(n9863) );
  ND2HHD U14243 ( .I1(n12995), .I2(n8264), .O(n13050) );
  ND2HHD U14244 ( .I1(n9866), .I2(n8305), .O(n6259) );
  ND2HHD U14245 ( .I1(n9383), .I2(n7723), .O(n10759) );
  ND2KHD U14246 ( .I1(n7032), .I2(n13442), .O(n9873) );
  INVCHD U14247 ( .I(n12431), .O(n9875) );
  NR2GHD U14248 ( .I1(n9876), .I2(n13192), .O(n13193) );
  ND2HHD U14249 ( .I1(n10080), .I2(n12376), .O(n9876) );
  ND3EHD U14250 ( .I1(n9879), .I2(n9880), .I3(n9881), .O(n9877) );
  ND2HHD U14251 ( .I1(n11584), .I2(_i_CLEFIA128_state_reg _1), .O(n9890) );
  NR2IHD U14252 ( .I1(n7674), .I2(n10471), .O(n11022) );
  OA13EHD U14253 ( .B1(n10272), .B2(n10273), .B3(n9899), .A1(n12462), .O(n10274) );
  ND3EHD U14254 ( .I1(n9908), .I2(n9907), .I3(n10560), .O(n9904) );
  ND2CHD U14255 ( .I1(n12239), .I2(n13004), .O(n9910) );
  XOR2HHD U14256 ( .I1(n13266), .I2(n13267), .O(n9913) );
  ND2HHD U14257 ( .I1(n12713), .I2(n9916), .O(n10902) );
  ND2KHD U14258 ( .I1(n7038), .I2(n6909), .O(n13005) );
  NR2IHD U14259 ( .I1(n8212), .I2(n10328), .O(n10644) );
  ND2KHD U14260 ( .I1(n7039), .I2(n8188), .O(n12730) );
  XNR2HHD U14261 ( .I1(DOUT_65), .I2(n9923), .O(n14228) );
  NR2GHD U14262 ( .I1(n10750), .I2(n9924), .O(n10751) );
  XOR2HHD U14263 ( .I1(n10158), .I2(n9930), .O(n13040) );
  ND2HHD U14264 ( .I1(n9934), .I2(n10165), .O(n9933) );
  ND2HHD U14265 ( .I1(n10882), .I2(n12788), .O(n9940) );
  ND2HHD U14266 ( .I1(n10305), .I2(_i_CLEFIA128_state_reg _1), .O(n9943) );
  AN3HHD U14267 ( .I1(n10452), .I2(n10939), .I3(n10090), .O(n12809) );
  ND2KHD U14268 ( .I1(n8797), .I2(_i_CLEFIA128_keyK _43), .O(n10157) );
  INVLHD U14269 ( .I(_i_CLEFIA128_keyL _107), .O(n14817) );
  ND2HHD U14270 ( .I1(n10323), .I2(_i_CLEFIA128_state_reg _1), .O(n9951) );
  OR3HHD U14271 ( .I1(n12849), .I2(n10830), .I3(n10829), .O(n9952) );
  XNR3EHD U14272 ( .I1(n9955), .I2(n14016), .I3(n12828), .O(n9954) );
  XOR2HHD U14273 ( .I1(n13911), .I2(n7256), .O(n9957) );
  ND2HHD U14274 ( .I1(n9966), .I2(n12474), .O(n9965) );
  ND2HHD U14275 ( .I1(n10629), .I2(n6807), .O(n9966) );
  XNR2HHD U14276 ( .I1(n9970), .I2(n14491), .O(n14492) );
  OR2EHD U14277 ( .I1(n8118), .I2(n9973), .O(n13364) );
  ND2HHD U14278 ( .I1(n9976), .I2(_i_CLEFIA128_state_reg _1), .O(n10118) );
  ND2HHD U14279 ( .I1(_i_CLEFIA128_keyK _11), .I2(n8797), .O(n9977) );
  INVLHD U14280 ( .I(_i_CLEFIA128_keyL _11), .O(n14939) );
  ND3EHD U14281 ( .I1(n9981), .I2(n8267), .I3(n12028), .O(n9980) );
  XOR2HHD U14282 ( .I1(n9985), .I2(n14344), .O(n10180) );
  ND2HHD U14283 ( .I1(n11864), .I2(n9988), .O(n9987) );
  INVCHD U14284 ( .I(n9995), .O(n9994) );
  ND2HHD U14285 ( .I1(n8202), .I2(n11226), .O(n10358) );
  ND2CHD U14286 ( .I1(n9747), .I2(n9998), .O(n13579) );
  XNR3EHD U14287 ( .I1(n10151), .I2(n10150), .I3(n7932), .O(n10000) );
  OR3HHD U14288 ( .I1(n11682), .I2(n12075), .I3(n11678), .O(n13810) );
  ND2HHD U14289 ( .I1(n12030), .I2(n8185), .O(n12934) );
  OR2EHD U14290 ( .I1(n13494), .I2(n10002), .O(n10297) );
  ND2HHD U14291 ( .I1(n10005), .I2(n6543), .O(n13129) );
  ND3EHD U14292 ( .I1(n13144), .I2(n12032), .I3(n10005), .O(n12033) );
  ND3EHD U14293 ( .I1(n9886), .I2(n13125), .I3(n10007), .O(n13617) );
  ND2HHD U14294 ( .I1(n10010), .I2(n14224), .O(n6153) );
  BUFQHD U14295 ( .I(n10791), .O(n10011) );
  ND3EHD U14296 ( .I1(n10016), .I2(n11263), .I3(n10015), .O(n10014) );
  ND2HHD U14297 ( .I1(n10775), .I2(n11221), .O(n10024) );
  XNR2HHD U14298 ( .I1(n10031), .I2(n10321), .O(n10030) );
  ND2KHD U14299 ( .I1(n10036), .I2(n6913), .O(n12305) );
  OAI12CHD U14300 ( .B1(n6790), .B2(n10279), .A1(n12474), .O(n10038) );
  ND2HHD U14301 ( .I1(n10040), .I2(n10041), .O(n6218) );
  AN2HHD U14302 ( .I1(n11400), .I2(n11399), .O(n10053) );
  ND2HHD U14303 ( .I1(n10061), .I2(n14153), .O(n6100) );
  MUX2HHD U14304 ( .A(n14146), .B(n14145), .S(n9836), .O(n10061) );
  ND3EHD U14305 ( .I1(n12559), .I2(n12765), .I3(n10073), .O(n10067) );
  ND2KHD U14306 ( .I1(n10057), .I2(n7014), .O(n11504) );
  INVCHD U14307 ( .I(DOUT_0), .O(n10075) );
  ND2KHD U14308 ( .I1(n10874), .I2(n10011), .O(n12538) );
  ND2HHD U14309 ( .I1(n10079), .I2(n10078), .O(n6115) );
  ND2HHD U14310 ( .I1(n10082), .I2(n10081), .O(n6106) );
  XOR2HHD U14311 ( .I1(n14244), .I2(n14246), .O(n10083) );
  ND2KHD U14312 ( .I1(n7398), .I2(n11049), .O(n12726) );
  ND2KHD U14313 ( .I1(n8904), .I2(n7039), .O(n11506) );
  XOR2HHD U14314 ( .I1(n14016), .I2(n14014), .O(n10086) );
  XNR2HHD U14315 ( .I1(n14013), .I2(n14017), .O(n10087) );
  ND2KHD U14316 ( .I1(n10202), .I2(n10200), .O(n10091) );
  ND3EHD U14317 ( .I1(n13457), .I2(n13430), .I3(n10094), .O(n10093) );
  AN2CHD U14318 ( .I1(n10745), .I2(n10219), .O(n10451) );
  OR3HHD U14319 ( .I1(n12441), .I2(n12242), .I3(n12243), .O(n13437) );
  ND2HHD U14320 ( .I1(n12235), .I2(n12989), .O(n10103) );
  ND2HHD U14321 ( .I1(n13018), .I2(n12989), .O(n12435) );
  ND2KHD U14322 ( .I1(n10599), .I2(n7671), .O(n12480) );
  ND2KHD U14323 ( .I1(n7671), .I2(n11274), .O(n11553) );
  OR3HHD U14324 ( .I1(n12919), .I2(n13124), .I3(n12918), .O(n13587) );
  ND2HHD U14325 ( .I1(n12127), .I2(n12291), .O(n12917) );
  ND3EHD U14326 ( .I1(n12740), .I2(n6891), .I3(n10518), .O(n11480) );
  ND2HHD U14327 ( .I1(n13018), .I2(n13459), .O(n12234) );
  OA13EHD U14328 ( .B1(n11538), .B2(n11537), .B3(n11536), .A1(n12462), .O(n11539) );
  ND2KHD U14329 ( .I1(n12327), .I2(n9676), .O(n13028) );
  ND3EHD U14330 ( .I1(n11019), .I2(n11380), .I3(n11379), .O(n12574) );
  ND2HHD U14331 ( .I1(n11018), .I2(n7398), .O(n11364) );
  MUX2HHD U14332 ( .A(n13793), .B(n13792), .S(n14525), .O(n13801) );
  ND2KHD U14333 ( .I1(n12129), .I2(n11995), .O(n13602) );
  OR3HHD U14334 ( .I1(n13656), .I2(n13655), .I3(n13654), .O(n13848) );
  ND3EHD U14335 ( .I1(n12027), .I2(n7031), .I3(n13629), .O(n13176) );
  NR2IHD U14336 ( .I1(n9857), .I2(n12000), .O(n12056) );
  OR3HHD U14337 ( .I1(n10697), .I2(n10698), .I3(n11311), .O(n10708) );
  XOR2HHD U14338 ( .I1(_i_CLEFIA128_keyL _104), .I2(n11869), .O(n11873) );
  ND2HHD U14339 ( .I1(n11360), .I2(n11333), .O(n11396) );
  OR3HHD U14340 ( .I1(n11020), .I2(n10484), .I3(n11504), .O(n10485) );
  ND2HHD U14341 ( .I1(n7900), .I2(n12456), .O(n11131) );
  ND2HHD U14342 ( .I1(n12944), .I2(n13608), .O(n13110) );
  XOR2HHD U14343 ( .I1(_i_CLEFIA128_CON_T_x _8), .I2(DOUT_104), .O(n11870));
  XOR2HHD U14344 ( .I1(n14103), .I2(n9013), .O(n14803) );
  ND2KHD U14345 ( .I1(n10318), .I2(n10668), .O(n12620) );
  ND3EHD U14346 ( .I1(n11037), .I2(n7115), .I3(n11036), .O(n11039) );
  NR2EHD U14347 ( .I1(n12218), .I2(n12435), .O(n13438) );
  ND2KHD U14348 ( .I1(n9903), .I2(n11274), .O(n10588) );
  ND2HHD U14349 ( .I1(n9676), .I2(n7032), .O(n12350) );
  MUX2HHD U14350 ( .A(n14232), .B(n14231), .S(n15054), .O(n14240) );
  MUX2HHD U14351 ( .A(n14390), .B(n14389), .S(n9540), .O(n14398) );
  ND3EHD U14352 ( .I1(n11625), .I2(n11626), .I3(n13083), .O(n11627) );
  ND2KHD U14353 ( .I1(n9684), .I2(n12829), .O(n10945) );
  ND2HHD U14354 ( .I1(n13367), .I2(n8357), .O(n10125) );
  ND2HHD U14355 ( .I1(n7830), .I2(n9676), .O(n13444) );
  OAI112BHD U14356 ( .C1(n12292), .C2(n10130), .A1(n6529), .B1(n13628), .O(n12295) );
  OR3HHD U14357 ( .I1(n13115), .I2(n13114), .I3(n10133), .O(n13116) );
  OR3HHD U14358 ( .I1(n12395), .I2(n10133), .I3(n12394), .O(n13173) );
  ND2HHD U14359 ( .I1(n12915), .I2(n9580), .O(n13627) );
  NR3BHD U14360 ( .I1(n12400), .I2(n12117), .I3(n10135), .O(n10134) );
  ND2HHD U14361 ( .I1(n12637), .I2(n12617), .O(n10137) );
  ND2HHD U14362 ( .I1(n10794), .I2(n12517), .O(n12617) );
  XNR2HHD U14363 ( .I1(DOUT_76), .I2(n8757), .O(n10147) );
  XOR2HHD U14364 ( .I1(n14328), .I2(n9923), .O(n10150) );
  ND2HHD U14365 ( .I1(n12912), .I2(n13585), .O(n13112) );
  XNR3EHD U14366 ( .I1(n7129), .I2(n10160), .I3(n10159), .O(n10158) );
  NR2GHD U14367 ( .I1(n13108), .I2(n12949), .O(n14996) );
  ND3EHD U14368 ( .I1(n10564), .I2(n10566), .I3(n10565), .O(n10163) );
  INVLHD U14369 ( .I(_i_CLEFIA128_keyL _81), .O(n15069) );
  ND2KHD U14370 ( .I1(n12424), .I2(n9430), .O(n13373) );
  ND2HHD U14371 ( .I1(n10247), .I2(n10316), .O(n10168) );
  ND2HHD U14372 ( .I1(n12736), .I2(n11512), .O(n12758) );
  ND3EHD U14373 ( .I1(n12120), .I2(n9207), .I3(n9456), .O(n10183) );
  ND2HHD U14374 ( .I1(n10192), .I2(n7005), .O(n6216) );
  ND2KHD U14375 ( .I1(n9801), .I2(n8180), .O(n11485) );
  ND2HHD U14376 ( .I1(n10123), .I2(n8215), .O(n12797) );
  ND2HHD U14377 ( .I1(n10219), .I2(n9684), .O(n12714) );
  ND2HHD U14378 ( .I1(n13442), .I2(n7830), .O(n12955) );
  OR3HHD U14379 ( .I1(n12336), .I2(n12337), .I3(n13029), .O(n10236) );
  OR3HHD U14380 ( .I1(n10237), .I2(n11280), .I3(n11279), .O(n12475) );
  NR2IHD U14381 ( .I1(n10593), .I2(n9733), .O(n10719) );
  OR3HHD U14382 ( .I1(n11392), .I2(n11393), .I3(n11391), .O(n11394) );
  INVCKGHD U14383 ( .I(n10553), .O(n10249) );
  ND2KHD U14384 ( .I1(n10712), .I2(n8179), .O(n10252) );
  XOR2HHD U14385 ( .I1(_i_CLEFIA128_keyL _92), .I2(n10258), .O(n10257) );
  ND2HHD U14386 ( .I1(_i_CLEFIA128_keyK _92), .I2(n8797), .O(n10258) );
  ND2HHD U14387 ( .I1(n11496), .I2(n11360), .O(n12724) );
  ND2HHD U14388 ( .I1(n7217), .I2(n7507), .O(n12623) );
  OR2EHD U14389 ( .I1(n11434), .I2(n12459), .O(n10273) );
  OAI12CHD U14390 ( .B1(n10278), .B2(n10276), .A1(n12491), .O(n10275) );
  ND3EHD U14391 ( .I1(n10280), .I2(n8335), .I3(n12467), .O(n10279) );
  AN2HHD U14392 ( .I1(n8413), .I2(n12466), .O(n10280) );
  ND2KHD U14393 ( .I1(n10123), .I2(n8916), .O(n10964) );
  XOR2HHD U14394 ( .I1(_i_CLEFIA128_keyL _91), .I2(n10289), .O(n10307) );
  ND2HHD U14395 ( .I1(_i_CLEFIA128_keyK _91), .I2(n8797), .O(n10289) );
  ND2KHD U14396 ( .I1(n11176), .I2(n11274), .O(n11284) );
  XOR2HHD U14397 ( .I1(n14171), .I2(n14029), .O(n14030) );
  ND2KHD U14398 ( .I1(n8214), .I2(n9430), .O(n13018) );
  OA13EHD U14399 ( .B1(n13588), .B2(n13586), .B3(n13587), .A1(n13585), .O(n13611) );
  NR2GHD U14400 ( .I1(n11653), .I2(n11652), .O(n14065) );
  ND2HHD U14401 ( .I1(n12980), .I2(n13458), .O(n13051) );
  ND2KHD U14402 ( .I1(n8210), .I2(n7292), .O(n14070) );
  ND2HHD U14403 ( .I1(n12902), .I2(n12291), .O(n12401) );
  ND2KHD U14404 ( .I1(n10794), .I2(n9659), .O(n11233) );
  INVMHD U14405 ( .I(_i_CLEFIA128_keyL _43), .O(n15191) );
  ND2HHD U14406 ( .I1(n8183), .I2(n12291), .O(n13128) );
  XNR2KHD U14407 ( .I1(n14493), .I2(n14492), .O(n15486) );
  ND2HHD U14408 ( .I1(n8196), .I2(n8178), .O(n12306) );
  ND2KHD U14409 ( .I1(n12129), .I2(n12915), .O(n12268) );
  ND2KHD U14410 ( .I1(n11049), .I2(n9801), .O(n12564) );
  XNR2HHD U14411 ( .I1(n14143), .I2(n13702), .O(n14615) );
  XNR2KHD U14412 ( .I1(n10398), .I2(n10397), .O(n12864) );
  ND2KHD U14413 ( .I1(n11948), .I2(n7032), .O(n13366) );
  ND2KHD U14414 ( .I1(n11948), .I2(n12251), .O(n13398) );
  ND2KHD U14415 ( .I1(n11948), .I2(n12226), .O(n13021) );
  AN2KHD U14416 ( .I1(n6803), .I2(n11245), .O(n12646) );
  AN2KHD U14417 ( .I1(n12335), .I2(n12349), .O(n13431) );
  INVMHD U14418 ( .I(_i_CLEFIA128_keyL _68), .O(n14931) );
  ND2KHD U14419 ( .I1(n7038), .I2(n7032), .O(n13447) );
  NR2IHD U14420 ( .I1(n9992), .I2(n10429), .O(n12836) );
  ND2KHD U14421 ( .I1(n10095), .I2(n12127), .O(n12935) );
  NR2GHD U14422 ( .I1(n10779), .I2(n11259), .O(n12650) );
  ND2KHD U14423 ( .I1(n11681), .I2(n8178), .O(n12302) );
  ND2KHD U14424 ( .I1(n12127), .I2(n12915), .O(n13122) );
  AN2KHD U14425 ( .I1(n12324), .I2(n12349), .O(n13458) );
  ND2KHD U14426 ( .I1(n13132), .I2(n11995), .O(n13187) );
  ND2HHD U14427 ( .I1(n12123), .I2(n13613), .O(n12260) );
  NR2GHD U14428 ( .I1(n12234), .I2(n12233), .O(n12418) );
  NR2EHD U14429 ( .I1(n10131), .I2(n9777), .O(n12930) );
  ND2KHD U14430 ( .I1(n12125), .I2(n13132), .O(n13194) );
  ND2KHD U14431 ( .I1(n11274), .I2(n12484), .O(n11438) );
  ND2KHD U14432 ( .I1(n9964), .I2(n12484), .O(n11552) );
  ND2KHD U14433 ( .I1(n12383), .I2(n10095), .O(n13590) );
  ND2HHD U14434 ( .I1(n9694), .I2(n9050), .O(n11337) );
  ND2HHD U14435 ( .I1(n13573), .I2(n12945), .O(n13618) );
  ND2KHD U14436 ( .I1(n12900), .I2(n8185), .O(n13573) );
  ND2HHD U14437 ( .I1(n12423), .I2(n12251), .O(n12436) );
  ND3EHD U14438 ( .I1(n10596), .I2(n10598), .I3(n10597), .O(n11310) );
  ND2KHD U14439 ( .I1(n9628), .I2(n8210), .O(n14081) );
  ND2KHD U14440 ( .I1(n11906), .I2(n12251), .O(n13439) );
  ND2KHD U14441 ( .I1(n12498), .I2(n8767), .O(n12502) );
  ND2KHD U14442 ( .I1(n9699), .I2(n12902), .O(n13589) );
  ND2HHD U14443 ( .I1(n9626), .I2(n10973), .O(n10990) );
  ND2KHD U14444 ( .I1(n12900), .I2(n12129), .O(n13613) );
  ND2KHD U14445 ( .I1(n10599), .I2(n10600), .O(n11531) );
  ND2KHD U14446 ( .I1(n9559), .I2(n8191), .O(n10966) );
  NR2GHD U14447 ( .I1(n10803), .I2(n6839), .O(n10669) );
  ND2KHD U14448 ( .I1(n11176), .I2(n6873), .O(n11292) );
  ND2KHD U14449 ( .I1(n12561), .I2(n9050), .O(n12731) );
  ND2KHD U14450 ( .I1(n7161), .I2(n9659), .O(n12621) );
  AN2HHD U14451 ( .I1(n11454), .I2(n11455), .O(n12467) );
  ND2HHD U14452 ( .I1(n12038), .I2(n12037), .O(n12941) );
  NR2EHD U14453 ( .I1(n12036), .I2(n12035), .O(n12037) );
  ND2KHD U14454 ( .I1(n12129), .I2(n12030), .O(n12945) );
  ND2KHD U14455 ( .I1(n10973), .I2(n9800), .O(n11178) );
  ND2KHD U14456 ( .I1(n11766), .I2(n8210), .O(n13084) );
  ND2KHD U14457 ( .I1(n12900), .I2(n12902), .O(n13628) );
  ND2KHD U14458 ( .I1(n8214), .I2(n7032), .O(n13448) );
  ND2KHD U14459 ( .I1(n7039), .I2(n11335), .O(n12577) );
  INVGHD U14460 ( .I(n9186), .O(n11764) );
  ND2HHD U14461 ( .I1(n9186), .I2(n9184), .O(n13223) );
  ND2HHD U14462 ( .I1(n9186), .I2(n11818), .O(n14052) );
  ND2KHD U14463 ( .I1(n7034), .I2(n9186), .O(n13099) );
  ND2KHD U14464 ( .I1(n12423), .I2(n12226), .O(n13372) );
  ND2HHD U14465 ( .I1(n11679), .I2(n6831), .O(n11682) );
  ND2KHD U14466 ( .I1(n11713), .I2(n8178), .O(n13510) );
  ND2KHD U14467 ( .I1(n7398), .I2(n7039), .O(n11510) );
  ND2KHD U14468 ( .I1(n12902), .I2(n11995), .O(n13125) );
  ND2KHD U14469 ( .I1(n10802), .I2(n10668), .O(n10783) );
  ND2KHD U14470 ( .I1(n10600), .I2(n11274), .O(n11459) );
  ND2KHD U14471 ( .I1(n11681), .I2(n9807), .O(n13838) );
  ND2KHD U14472 ( .I1(n12561), .I2(n9898), .O(n12737) );
  ND2KHD U14473 ( .I1(n7039), .I2(n9801), .O(n12586) );
  ND2KHD U14474 ( .I1(n10318), .I2(n9659), .O(n12537) );
  ND2KHD U14475 ( .I1(n9807), .I2(n13521), .O(n12309) );
  ND2KHD U14476 ( .I1(n8180), .I2(n7398), .O(n12766) );
  ND2KHD U14477 ( .I1(n9897), .I2(n8188), .O(n12559) );
  ND2KHD U14478 ( .I1(n8209), .I2(n12145), .O(n13681) );
  ND2KHD U14479 ( .I1(n8183), .I2(n10095), .O(n13592) );
  ND2KHD U14480 ( .I1(n8183), .I2(n12030), .O(n13591) );
  AO22CHD U14481 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _114), .B1(n15504), .B2(_i_CLEFIA128_keyK _50), .O(n10292) );
  AN2EHD U14482 ( .I1(n13399), .I2(n13398), .O(n13402) );
  INVJHD U14483 ( .I(_i_CLEFIA128_keyL _60), .O(n14936) );
  ND2DHD U14484 ( .I1(n15336), .I2(n15324), .O(n15334) );
  NR2GHD U14485 ( .I1(_i_CLEFIA128_rndcnt_reg _3), .I2(_i_CLEFIA128_rndcnt_reg _2), .O(n14419) );
  AN2HHD U14486 ( .I1(n14419), .I2(n10298), .O(n13278) );
  NR2IHD U14487 ( .I1(n7389), .I2(n13287), .O(n14688) );
  ND2HHD U14488 ( .I1(n10301), .I2(_i_CLEFIA128_state_reg _1), .O(n14685) );
  ND2KHD U14489 ( .I1(_i_CLEFIA128_rndcnt_reg _0), .I2(n8797), .O(n11979) );
  BUFQHD U14490 ( .I(n11979), .O(n14707) );
  XNR2EHD U14491 ( .I1(_i_CLEFIA128_CON_T_xi _11), .I2(DOUT_60), .O(n10312));
  ND2DHD U14492 ( .I1(_i_CLEFIA128_keyK _26), .I2(_i_CLEFIA128_keyL _26), .O(n10320) );
  ND2DHD U14493 ( .I1(n10798), .I2(n12609), .O(n10331) );
  INVDHD U14494 ( .I(n10328), .O(n12638) );
  ND2DHD U14495 ( .I1(n7507), .I2(n12638), .O(n10329) );
  INVDHD U14496 ( .I(n10332), .O(n10632) );
  INVDHD U14497 ( .I(_i_CLEFIA128_keyK _30), .O(n13909) );
  NR2CHD U14498 ( .I1(n13909), .I2(n14707), .O(n10339) );
  XNR2KHD U14499 ( .I1(n10343), .I2(n10342), .O(n11216) );
  XOR2EHD U14500 ( .I1(_i_CLEFIA128_CON_T_x _0), .I2(DOUT_63), .O(n10353) );
  INVDHD U14501 ( .I(_i_CLEFIA128_keyK _31), .O(n13790) );
  MXL2CHD U14502 ( .A(n10349), .B(n10348), .S(_i_CLEFIA128_keyL _31), .OB(n10350) );
  XNR2KHD U14503 ( .I1(n10353), .I2(n10352), .O(n11230) );
  INVDHD U14504 ( .I(n10363), .O(n10773) );
  ND2DHD U14505 ( .I1(n10773), .I2(n10668), .O(n10364) );
  NR2CHD U14506 ( .I1(n10365), .I2(n12653), .O(n10366) );
  NR3BHD U14507 ( .I1(n6846), .I2(n10801), .I3(n10370), .O(n10374) );
  ND2DHD U14508 ( .I1(n11063), .I2(n10851), .O(n10372) );
  NR2CHD U14509 ( .I1(n10372), .I2(n10371), .O(n10373) );
  NR2CHD U14510 ( .I1(n10375), .I2(n10801), .O(n10376) );
  ND2DHD U14511 ( .I1(n12619), .I2(n11070), .O(n10377) );
  INVDHD U14512 ( .I(n10859), .O(n10387) );
  NR3BHD U14513 ( .I1(n6906), .I2(n10387), .I3(n12626), .O(n10388) );
  XOR2EHD U14514 ( .I1(_i_CLEFIA128_CON_T_x _7), .I2(DOUT_46), .O(n10398) );
  INVDHD U14515 ( .I(_i_CLEFIA128_keyK _14), .O(n13949) );
  MXL2CHD U14516 ( .A(n10394), .B(n10393), .S(_i_CLEFIA128_keyL _14), .OB(n10395) );
  INVDHD U14517 ( .I(_i_CLEFIA128_keyK _15), .O(n14784) );
  NR2CHD U14518 ( .I1(n10422), .I2(n12780), .O(n10423) );
  NR2CHD U14519 ( .I1(n10820), .I2(n12799), .O(n10434) );
  INVDHD U14520 ( .I(n10964), .O(n10430) );
  NR2CHD U14521 ( .I1(n12836), .I2(n10430), .O(n10433) );
  NR2CHD U14522 ( .I1(n12808), .I2(n8915), .O(n10432) );
  ND2DHD U14523 ( .I1(n6879), .I2(n9844), .O(n10443) );
  ND2DHD U14524 ( .I1(n10939), .I2(n10123), .O(n10958) );
  ND2DHD U14525 ( .I1(n12829), .I2(n10939), .O(n10961) );
  ND2DHD U14526 ( .I1(n12856), .I2(n12717), .O(n12685) );
  INVDHD U14527 ( .I(n12689), .O(n10447) );
  INVDHD U14528 ( .I(n6767), .O(n10745) );
  XOR2EHD U14529 ( .I1(_i_CLEFIA128_CON_T_x _12), .I2(DOUT_35), .O(n10455));
  XNR2EHD U14530 ( .I1(_i_CLEFIA128_CON_T_x _14), .I2(DOUT_37), .O(n10460));
  NR2CHD U14531 ( .I1(n12552), .I2(n10475), .O(n10478) );
  ND2DHD U14532 ( .I1(n12578), .I2(n11485), .O(n10476) );
  ND3CHD U14533 ( .I1(n8463), .I2(n10478), .I3(n10477), .O(n10506) );
  ND2DHD U14534 ( .I1(n7146), .I2(n11340), .O(n10482) );
  ND3CHD U14535 ( .I1(n11322), .I2(n11484), .I3(n11100), .O(n10505) );
  NR2CHD U14536 ( .I1(n11488), .I2(n11033), .O(n10486) );
  ND2DHD U14537 ( .I1(n12556), .I2(n10486), .O(n10504) );
  XOR2EHD U14538 ( .I1(_i_CLEFIA128_CON_T_x _0), .I2(DOUT_39), .O(n10496) );
  OR2B1CHD U14539 ( .I1(_i_CLEFIA128_keyK _7), .B1(n8691), .O(n10490) );
  INVDHD U14540 ( .I(_i_CLEFIA128_keyK _7), .O(n14772) );
  MXL2CHD U14541 ( .A(n10492), .B(n10491), .S(_i_CLEFIA128_keyL _7), .OB(n10493) );
  XOR2EHD U14542 ( .I1(_i_CLEFIA128_CON_T_xi _13), .I2(DOUT_38), .O(n10503));
  INVDHD U14543 ( .I(_i_CLEFIA128_keyK _6), .O(n14011) );
  OAI13BHD U14544 ( .B1(n10506), .B2(n10505), .B3(n10504), .A1(n11500), .O(n10543) );
  NR2CHD U14545 ( .I1(n10509), .I2(n10508), .O(n10511) );
  INVDHD U14546 ( .I(n12724), .O(n10510) );
  NR2CHD U14547 ( .I1(n11480), .I2(n12573), .O(n10524) );
  INVDHD U14548 ( .I(n11504), .O(n11018) );
  ND2DHD U14549 ( .I1(n11378), .I2(n11335), .O(n10519) );
  AN3EHD U14550 ( .I1(n11410), .I2(n12747), .I3(n10519), .O(n10520) );
  ND3CHD U14551 ( .I1(n10535), .I2(n10520), .I3(n12726), .O(n10521) );
  NR2CHD U14552 ( .I1(n10521), .I2(n10522), .O(n10523) );
  ND2HHD U14553 ( .I1(n12731), .I2(n11333), .O(n12579) );
  ND3CHD U14554 ( .I1(n10533), .I2(n11506), .I3(n11358), .O(n10540) );
  OR3EHD U14555 ( .I1(n10540), .I2(n10539), .I3(n12761), .O(n10541) );
  INVMHD U14556 ( .I(_i_CLEFIA128_keyL _19), .O(n15263) );
  ND2HHD U14557 ( .I1(n10546), .I2(_i_CLEFIA128_state_reg _1), .O(n10547) );
  XOR2EHD U14558 ( .I1(_i_CLEFIA128_CON_T_reg_4 ), .I2(DOUT_52), .O(n10555));
  ND2KHD U14559 ( .I1(n8039), .I2(_i_CLEFIA128_keyK _20), .O(n10553) );
  XOR2EHD U14560 ( .I1(_i_CLEFIA128_CON_T_x _6), .I2(DOUT_53), .O(n10560) );
  OR2B1CHD U14561 ( .I1(n8797), .B1(_i_CLEFIA128_keyL _81), .O(n10565) );
  INVMHD U14562 ( .I(_i_CLEFIA128_keyL _17), .O(n14988) );
  ND2KHD U14563 ( .I1(n10973), .I2(n9964), .O(n12468) );
  INVDHD U14564 ( .I(_i_CLEFIA128_keyK _22), .O(n13984) );
  MXL2CHD U14565 ( .A(n10578), .B(n10577), .S(_i_CLEFIA128_keyL _22), .OB(n10579) );
  ND3CHD U14566 ( .I1(n12449), .I2(n12480), .I3(n9034), .O(n10584) );
  XOR2EHD U14567 ( .I1(_i_CLEFIA128_CON_T_x _8), .I2(DOUT_55), .O(n10610) );
  OR2B1CHD U14568 ( .I1(_i_CLEFIA128_keyK _23), .B1(n8691), .O(n10604) );
  INVDHD U14569 ( .I(_i_CLEFIA128_keyK _23), .O(n13881) );
  NR2CHD U14570 ( .I1(n13881), .I2(n7103), .O(n10605) );
  MXL2CHD U14571 ( .A(n10606), .B(n10605), .S(_i_CLEFIA128_keyL _23), .OB(n10607) );
  ND3CHD U14572 ( .I1(n10608), .I2(n10607), .I3(_i_CLEFIA128_state_reg _1), .O(n10609) );
  ND2DHD U14573 ( .I1(n11439), .I2(n9047), .O(n10612) );
  NR2CHD U14574 ( .I1(n12496), .I2(n10612), .O(n10614) );
  NR2CHD U14575 ( .I1(n11448), .I2(n8770), .O(n10613) );
  ND2DHD U14576 ( .I1(n10617), .I2(n9903), .O(n10618) );
  ND2DHD U14577 ( .I1(n11554), .I2(n11546), .O(n11179) );
  ND2DHD U14578 ( .I1(n8768), .I2(n10690), .O(n10624) );
  INVDHD U14579 ( .I(n11060), .O(n10635) );
  ND2DHD U14580 ( .I1(n10173), .I2(n7216), .O(n10637) );
  ND2DHD U14581 ( .I1(n10638), .I2(n12657), .O(n10640) );
  ND3CHD U14582 ( .I1(n9648), .I2(n10783), .I3(n11236), .O(n10642) );
  NR2CHD U14583 ( .I1(n10647), .I2(n11085), .O(n10648) );
  ND2DHD U14584 ( .I1(n10862), .I2(n6617), .O(n10652) );
  NR2CHD U14585 ( .I1(n10652), .I2(n10651), .O(n10653) );
  NR2CHD U14586 ( .I1(n10659), .I2(n10660), .O(n10661) );
  INVDHD U14587 ( .I(n11233), .O(n10666) );
  INVDHD U14588 ( .I(n10668), .O(n10670) );
  ND2DHD U14589 ( .I1(n6578), .I2(n7507), .O(n10672) );
  ND3CHD U14590 ( .I1(n10673), .I2(n11236), .I3(n10672), .O(n10675) );
  ND2DHD U14591 ( .I1(n12621), .I2(n12652), .O(n10674) );
  OR3HHD U14592 ( .I1(n12526), .I2(n10681), .I3(n10682), .O(n10684) );
  ND2DHD U14593 ( .I1(n10567), .I2(n10690), .O(n11520) );
  AN3EHD U14594 ( .I1(n11443), .I2(n6764), .I3(n11520), .O(n10691) );
  ND3CHD U14595 ( .I1(n10692), .I2(n10691), .I3(n12489), .O(n10693) );
  OA13EHD U14596 ( .B1(n10694), .B2(n10693), .B3(n11310), .A1(n12474), .O(n10710) );
  ND2DHD U14597 ( .I1(n8767), .I2(n11181), .O(n10699) );
  OAI12CHD U14598 ( .B1(n6567), .B2(n11183), .A1(n10699), .O(n10700) );
  AN2EHD U14599 ( .I1(n11312), .I2(n11318), .O(n12491) );
  AN2EHD U14600 ( .I1(n12456), .I2(n9034), .O(n10988) );
  ND3CHD U14601 ( .I1(n10717), .I2(n10716), .I3(n10715), .O(n10718) );
  NR2CHD U14602 ( .I1(n8179), .I2(n10720), .O(n12483) );
  ND2DHD U14603 ( .I1(n9903), .I2(n12483), .O(n11191) );
  ND2DHD U14604 ( .I1(n10746), .I2(n10745), .O(n10747) );
  NR2CHD U14605 ( .I1(n10749), .I2(n10748), .O(n10752) );
  ND3CHD U14606 ( .I1(n8423), .I2(n8812), .I3(n6706), .O(n10765) );
  INVDHD U14607 ( .I(n10760), .O(n10762) );
  NR2CHD U14608 ( .I1(n9561), .I2(n7216), .O(n10793) );
  NR2CHD U14609 ( .I1(n10795), .I2(n11065), .O(n10873) );
  ND3CHD U14610 ( .I1(n12878), .I2(n12864), .I3(n10825), .O(n10809) );
  NR2CHD U14611 ( .I1(n12789), .I2(n12675), .O(n10817) );
  ND2DHD U14612 ( .I1(n8812), .I2(n12864), .O(n10830) );
  ND3CHD U14613 ( .I1(n11221), .I2(n12538), .I3(n11216), .O(n10834) );
  NR3BHD U14614 ( .I1(n10834), .I2(n12529), .I3(n12658), .O(n10841) );
  ND3CHD U14615 ( .I1(n10839), .I2(n10840), .I3(n10841), .O(n10854) );
  NR2CHD U14616 ( .I1(n10856), .I2(n10857), .O(n10858) );
  INVDHD U14617 ( .I(n10862), .O(n10865) );
  ND3CHD U14618 ( .I1(n11236), .I2(n6803), .I3(n9648), .O(n10864) );
  NR2CHD U14619 ( .I1(n10871), .I2(n10870), .O(n10872) );
  ND2DHD U14620 ( .I1(n10874), .I2(n12638), .O(n10875) );
  INVGHD U14621 ( .I(DATASET), .O(n10908) );
  NR2GHD U14622 ( .I1(MODE_0), .I2(n10908), .O(n10915) );
  ND2HHD U14623 ( .I1(n10915), .I2(n10909), .O(n10910) );
  NR2IHD U14624 ( .I1(n10910), .I2(BSY), .O(n12895) );
  NR2IHD U14625 ( .I1(MODE_1), .I2(BSY), .O(n10916) );
  AN2KHD U14626 ( .I1(n12895), .I2(ENCDEC), .O(n13292) );
  AOI22BHD U14627 ( .A1(n7017), .A2(KEY_4), .B1(n13292), .B2(n10918), .O(n10919) );
  OAI112BHD U14628 ( .C1(n10912), .C2(n10921), .A1(n10920), .B1(n10919), .O(n10926) );
  OAI22CHD U14629 ( .A1(n14814), .A2(n15450), .B1(n15512), .B2(n14983), .O(n10925) );
  BUFQHD U14630 ( .I(n15450), .O(n15513) );
  AOI22BHD U14631 ( .A1(n7017), .A2(KEY_20), .B1(n13292), .B2(n10929), .O(n10930) );
  NR2CHD U14632 ( .I1(n9991), .I2(n10938), .O(n12709) );
  AN2EHD U14633 ( .I1(n10939), .I2(n8191), .O(n10940) );
  NR2CHD U14634 ( .I1(n12709), .I2(n10940), .O(n10941) );
  ND3CHD U14635 ( .I1(n10941), .I2(n6643), .I3(n12710), .O(n10942) );
  ND2DHD U14636 ( .I1(n9003), .I2(n8236), .O(n10944) );
  ND2DHD U14637 ( .I1(n8508), .I2(n12866), .O(n10949) );
  NR3BHD U14638 ( .I1(n10950), .I2(n10949), .I3(n10948), .O(n10955) );
  NR2CHD U14639 ( .I1(n12799), .I2(n10952), .O(n10953) );
  INVDHD U14640 ( .I(n12714), .O(n10956) );
  NR3BHD U14641 ( .I1(n12836), .I2(n10957), .I3(n10956), .O(n10968) );
  ND3CHD U14642 ( .I1(n10981), .I2(n10982), .I3(n10983), .O(n10984) );
  INVDHD U14643 ( .I(n11546), .O(n10995) );
  NR2CHD U14644 ( .I1(n10995), .I2(n12457), .O(n10999) );
  NR2CHD U14645 ( .I1(n10997), .I2(n10996), .O(n10998) );
  NR3BHD U14646 ( .I1(n11159), .I2(n11001), .I3(n11305), .O(n11003) );
  NR2CHD U14647 ( .I1(n11432), .I2(n11193), .O(n11002) );
  NR2CHD U14648 ( .I1(n11007), .I2(n11160), .O(n11011) );
  NR2CHD U14649 ( .I1(n11009), .I2(n11008), .O(n11010) );
  ND2DHD U14650 ( .I1(n11049), .I2(n11336), .O(n11014) );
  ND2KHD U14651 ( .I1(n11349), .I2(n10073), .O(n11401) );
  ND2DHD U14652 ( .I1(n11049), .I2(n6895), .O(n11023) );
  INVDHD U14653 ( .I(n9750), .O(n11048) );
  ND2DHD U14654 ( .I1(n9897), .I2(n11048), .O(n12566) );
  AN2EHD U14655 ( .I1(n12747), .I2(n12752), .O(n11479) );
  INVDHD U14656 ( .I(n11335), .O(n11030) );
  AN2EHD U14657 ( .I1(n12778), .I2(n12752), .O(n12591) );
  NR2CHD U14658 ( .I1(n11035), .I2(n11034), .O(n11036) );
  ND2DHD U14659 ( .I1(n11360), .I2(n11506), .O(n11041) );
  NR2CHD U14660 ( .I1(n11040), .I2(n11041), .O(n11042) );
  ND3CHD U14661 ( .I1(n12722), .I2(n11119), .I3(n11047), .O(n11056) );
  ND2DHD U14662 ( .I1(n11049), .I2(n11048), .O(n11507) );
  ND2DHD U14663 ( .I1(n11411), .I2(n11507), .O(n11050) );
  ND2DHD U14664 ( .I1(n12577), .I2(n11333), .O(n11053) );
  ND2DHD U14665 ( .I1(n11506), .I2(n12731), .O(n11052) );
  NR2CHD U14666 ( .I1(n11053), .I2(n11052), .O(n11054) );
  ND2DHD U14667 ( .I1(n12655), .I2(n12609), .O(n11061) );
  INVDHD U14668 ( .I(n11065), .O(n11067) );
  INVDHD U14669 ( .I(n11094), .O(n12751) );
  ND2DHD U14670 ( .I1(n12751), .I2(n7398), .O(n11096) );
  NR2GHD U14671 ( .I1(n9036), .I2(n11383), .O(n11099) );
  ND2DHD U14672 ( .I1(n11358), .I2(n12559), .O(n11104) );
  ND2DHD U14673 ( .I1(n12553), .I2(n8607), .O(n11103) );
  NR2CHD U14674 ( .I1(n11104), .I2(n11103), .O(n11105) );
  NR2CHD U14675 ( .I1(n11110), .I2(n11474), .O(n11113) );
  INVDHD U14676 ( .I(n11111), .O(n11112) );
  ND2DHD U14677 ( .I1(n7039), .I2(n11336), .O(n11120) );
  ND2DHD U14678 ( .I1(n11340), .I2(n11120), .O(n11122) );
  NR2CHD U14679 ( .I1(n11122), .I2(n11121), .O(n11123) );
  NR2CHD U14680 ( .I1(n11149), .I2(n11148), .O(n11150) );
  ND3CHD U14681 ( .I1(n7002), .I2(n11151), .I3(n11150), .O(n11152) );
  OA13EHD U14682 ( .B1(n11152), .B2(n11153), .B3(n11544), .A1(n12462), .O(n11154) );
  OA112EHD U14683 ( .C1(n11183), .C2(n11285), .A1(n12502), .B1(n11459), .O(n11167) );
  ND2DHD U14684 ( .I1(n11167), .I2(n8426), .O(n11172) );
  ND2DHD U14685 ( .I1(n6764), .I2(n12468), .O(n11170) );
  OR3EHD U14686 ( .I1(n11170), .I2(n11168), .I3(n11169), .O(n11171) );
  NR2CHD U14687 ( .I1(n11172), .I2(n11171), .O(n11173) );
  ND2DHD U14688 ( .I1(n11439), .I2(n11178), .O(n11180) );
  NR2CHD U14689 ( .I1(n11180), .I2(n11179), .O(n11185) );
  NR2CHD U14690 ( .I1(n11461), .I2(n11186), .O(n11198) );
  ND3CHD U14691 ( .I1(n11188), .I2(n11531), .I3(n12451), .O(n11189) );
  ND2DHD U14692 ( .I1(n11192), .I2(n11191), .O(n11194) );
  NR3BHD U14693 ( .I1(n11194), .I2(n11193), .I3(n11447), .O(n11196) );
  INVDHD U14694 ( .I(n12491), .O(n11195) );
  AO13EHD U14695 ( .B1(n11198), .B2(n11197), .B3(n11196), .A1(n11195), .O(n11199) );
  INVDHD U14696 ( .I(n11204), .O(n11208) );
  INVDHD U14697 ( .I(n11205), .O(n11206) );
  NR2CHD U14698 ( .I1(n11208), .I2(n11207), .O(n11209) );
  AN3EHD U14699 ( .I1(n11250), .I2(n11221), .I3(n12640), .O(n11213) );
  ND3CHD U14700 ( .I1(n12537), .I2(n9709), .I3(n11216), .O(n11218) );
  AN2EHD U14701 ( .I1(n12538), .I2(n12640), .O(n11227) );
  ND2DHD U14702 ( .I1(n12655), .I2(n11233), .O(n11239) );
  ND3CHD U14703 ( .I1(n11244), .I2(n12596), .I3(n11243), .O(n11246) );
  INVDHD U14704 ( .I(n11274), .O(n11275) );
  NR2CHD U14705 ( .I1(n11424), .I2(n11276), .O(n11277) );
  INVDHD U14706 ( .I(n8768), .O(n11286) );
  OA112EHD U14707 ( .C1(n11286), .C2(n11285), .A1(n11284), .B1(n9034), .O(n11288) );
  NR2CHD U14708 ( .I1(n11302), .I2(n11301), .O(n11303) );
  OR3EHD U14709 ( .I1(n11310), .I2(n11536), .I3(n11309), .O(n11320) );
  AN2B1CHD U14710 ( .I1(n11464), .B1(n11311), .O(n11317) );
  ND3CHD U14711 ( .I1(n11553), .I2(n9047), .I3(n11312), .O(n11313) );
  ND2DHD U14712 ( .I1(n11326), .I2(n11376), .O(n11327) );
  ND2DHD U14713 ( .I1(n12726), .I2(n12585), .O(n11331) );
  ND3CHD U14714 ( .I1(n12749), .I2(n12778), .I3(n11511), .O(n11330) );
  ND2DHD U14715 ( .I1(n11349), .I2(n11506), .O(n11338) );
  INVDHD U14716 ( .I(n11362), .O(n11343) );
  INVDHD U14717 ( .I(n11476), .O(n11347) );
  INVDHD U14718 ( .I(n11471), .O(n11346) );
  OA13EHD U14719 ( .B1(n11357), .B2(n11356), .B3(n11355), .A1(n12575), .O(n11363) );
  AN3EHD U14720 ( .I1(n9625), .I2(n11365), .I3(n11364), .O(n11366) );
  AN2EHD U14721 ( .I1(n12586), .I2(n11496), .O(n11370) );
  AN2EHD U14722 ( .I1(n12731), .I2(n11368), .O(n11369) );
  ND3CHD U14723 ( .I1(n11371), .I2(n11370), .I3(n11369), .O(n11372) );
  AN2HHD U14724 ( .I1(n11375), .I2(n12591), .O(n11390) );
  ND3CHD U14725 ( .I1(n11385), .I2(n11386), .I3(n9619), .O(n11387) );
  NR2CHD U14726 ( .I1(n11396), .I2(n11397), .O(n11400) );
  NR2CHD U14727 ( .I1(n11398), .I2(n12744), .O(n11399) );
  ND3CHD U14728 ( .I1(n12502), .I2(n11438), .I3(n11552), .O(n11423) );
  ND2DHD U14729 ( .I1(n8767), .I2(n8216), .O(n11430) );
  ND2DHD U14730 ( .I1(n6766), .I2(n6675), .O(n11437) );
  ND3CHD U14731 ( .I1(n11439), .I2(n11438), .I3(n11437), .O(n11441) );
  NR2CHD U14732 ( .I1(n11444), .I2(n11445), .O(n11446) );
  NR2CHD U14733 ( .I1(n11452), .I2(n8770), .O(n11455) );
  ND3CHD U14734 ( .I1(n11460), .I2(n12454), .I3(n12450), .O(n11462) );
  INVDHD U14735 ( .I(n12494), .O(n11465) );
  ND3CHD U14736 ( .I1(n11465), .I2(n11464), .I3(n11463), .O(n11466) );
  INVDHD U14737 ( .I(n12743), .O(n11473) );
  ND2DHD U14738 ( .I1(n6817), .I2(n12729), .O(n11486) );
  ND3CHD U14739 ( .I1(n12769), .I2(n6867), .I3(n11510), .O(n11516) );
  NR3BHD U14740 ( .I1(n11551), .I2(n11550), .I3(n11549), .O(n11558) );
  XOR2EHD U14741 ( .I1(_i_CLEFIA128_CON_T_x _14), .I2(DOUT_125), .O(n11566));
  XNR2KHD U14742 ( .I1(n11566), .I2(n11565), .O(n11647) );
  ND2DHD U14743 ( .I1(_i_CLEFIA128_keyK _57), .I2(_i_CLEFIA128_keyL _57), .O(n11567) );
  ND2KHD U14744 ( .I1(n8797), .I2(_i_CLEFIA128_keyK _122), .O(n11573) );
  XNR2EHD U14745 ( .I1(_i_CLEFIA128_CON_T_x _12), .I2(DOUT_123), .O(n11583));
  OR2B1CHD U14746 ( .I1(n8797), .B1(_i_CLEFIA128_keyL _123), .O(n11577) );
  XNR2KHD U14747 ( .I1(n11583), .I2(n11582), .O(n11612) );
  XOR2EHD U14748 ( .I1(_i_CLEFIA128_CON_T_x _0), .I2(DOUT_127), .O(n11601));
  INVDHD U14749 ( .I(_i_CLEFIA128_keyK _63), .O(n14754) );
  INVDHD U14750 ( .I(_i_CLEFIA128_keyK _62), .O(n13570) );
  NR2CHD U14751 ( .I1(n13570), .I2(n14707), .O(n11606) );
  MXL2CHD U14752 ( .A(n11607), .B(n11606), .S(_i_CLEFIA128_keyL _62), .OB(n11608) );
  ND3CHD U14753 ( .I1(n13469), .I2(n14049), .I3(n14052), .O(n11610) );
  NR2CHD U14754 ( .I1(n12202), .I2(n11610), .O(n11611) );
  ND3CHD U14755 ( .I1(n11822), .I2(n11611), .I3(n13229), .O(n11639) );
  INVDHD U14756 ( .I(n13099), .O(n11620) );
  ND2DHD U14757 ( .I1(n9597), .I2(n13100), .O(n11617) );
  ND3CHD U14758 ( .I1(n11764), .I2(n11628), .I3(n9184), .O(n11629) );
  ND2DHD U14759 ( .I1(n13096), .I2(n13083), .O(n11643) );
  ND3CHD U14760 ( .I1(n11645), .I2(n11822), .I3(n14047), .O(n11659) );
  INVDHD U14761 ( .I(n13096), .O(n11653) );
  XNR2EHD U14762 ( .I1(_i_CLEFIA128_CON_T_reg_4 ), .I2(DOUT_116), .O(n11660));
  XOR2EHD U14763 ( .I1(_i_CLEFIA128_CON_T_x _6), .I2(DOUT_117), .O(n11664));
  ND2DHD U14764 ( .I1(_i_CLEFIA128_keyK _51), .I2(_i_CLEFIA128_keyL _51), .O(n11666) );
  ND2DHD U14765 ( .I1(n8797), .I2(_i_CLEFIA128_keyK _51), .O(n11665) );
  ND3CHD U14766 ( .I1(n8310), .I2(n11675), .I3(n7389), .O(n11676) );
  INVDHD U14767 ( .I(_i_CLEFIA128_keyK _55), .O(n13765) );
  MXL2CHD U14768 ( .A(n11691), .B(n11690), .S(_i_CLEFIA128_keyL _55), .OB(n11692) );
  ND3CHD U14769 ( .I1(n11693), .I2(n11692), .I3(_i_CLEFIA128_state_reg _1), .O(n11694) );
  XOR2EHD U14770 ( .I1(_i_CLEFIA128_CON_T_x _7), .I2(DOUT_118), .O(n11705));
  INVDHD U14771 ( .I(_i_CLEFIA128_keyK _54), .O(n13995) );
  MXL2CHD U14772 ( .A(n11701), .B(n11700), .S(_i_CLEFIA128_keyL _54), .OB(n11702) );
  INVDHD U14773 ( .I(n11736), .O(n11727) );
  ND2DHD U14774 ( .I1(n13513), .I2(n11787), .O(n13647) );
  ND2DHD U14775 ( .I1(n9621), .I2(n13810), .O(n11734) );
  AN2EHD U14776 ( .I1(n11739), .I2(n6632), .O(n11740) );
  NR2CHD U14777 ( .I1(n13489), .I2(n11741), .O(n11742) );
  ND2DHD U14778 ( .I1(n14056), .I2(n14072), .O(n11746) );
  ND2DHD U14779 ( .I1(n9628), .I2(n13100), .O(n11747) );
  ND2DHD U14780 ( .I1(n13076), .I2(n13066), .O(n11748) );
  ND3CHD U14781 ( .I1(n13066), .I2(n8197), .I3(n14052), .O(n12205) );
  AN3EHD U14782 ( .I1(n13479), .I2(n14072), .I3(n13251), .O(n11759) );
  ND2DHD U14783 ( .I1(n11759), .I2(n11758), .O(n11760) );
  NR2CHD U14784 ( .I1(n12205), .I2(n11760), .O(n11765) );
  INVDHD U14785 ( .I(n11762), .O(n14060) );
  ND2HHD U14786 ( .I1(n11820), .I2(n13084), .O(n11829) );
  INVDHD U14787 ( .I(n11829), .O(n11769) );
  ND2DHD U14788 ( .I1(n9604), .I2(n7809), .O(n13812) );
  INVDHD U14789 ( .I(n13671), .O(n11788) );
  ND2DHD U14790 ( .I1(n13513), .I2(n13510), .O(n11790) );
  INVDHD U14791 ( .I(n11793), .O(n12171) );
  ND2DHD U14792 ( .I1(n7809), .I2(n12171), .O(n12069) );
  ND2DHD U14793 ( .I1(n6872), .I2(n7538), .O(n11795) );
  INVDHD U14794 ( .I(n8771), .O(n12159) );
  ND2DHD U14795 ( .I1(n7538), .I2(n9811), .O(n11806) );
  INVDHD U14796 ( .I(n6785), .O(n11812) );
  ND2DHD U14797 ( .I1(n8178), .I2(n7773), .O(n11816) );
  AN2EHD U14798 ( .I1(n14060), .I2(n11818), .O(n11819) );
  NR3BHD U14799 ( .I1(n13489), .I2(n11825), .I3(n11826), .O(n11828) );
  AN2EHD U14800 ( .I1(n13479), .I2(n13096), .O(n11827) );
  INVDHD U14801 ( .I(n13487), .O(n11830) );
  INVDHD U14802 ( .I(n11832), .O(n11833) );
  INVDHD U14803 ( .I(n11839), .O(n13231) );
  ND2DHD U14804 ( .I1(n13231), .I2(n9597), .O(n11842) );
  INVDHD U14805 ( .I(n13224), .O(n13483) );
  ND2DHD U14806 ( .I1(n13487), .I2(n14055), .O(n11847) );
  NR3BHD U14807 ( .I1(n13232), .I2(n13254), .I3(n11849), .O(n11850) );
  OA13EHD U14808 ( .B1(n11853), .B2(n13247), .B3(n13495), .A1(n14067), .O(n11854) );
  XNR2EHD U14809 ( .I1(_i_CLEFIA128_CON_T_xi _9), .I2(DOUT_107), .O(n11860));
  ND2DHD U14810 ( .I1(_i_CLEFIA128_keyK _40), .I2(_i_CLEFIA128_keyL _40), .O(n11868) );
  OAI112BHD U14811 ( .C1(n14707), .C2(n11868), .A1(n11867), .B1(_i_CLEFIA128_state_reg _1), .O(n11866) );
  XOR2EHD U14812 ( .I1(_i_CLEFIA128_CON_T_x _9), .I2(DOUT_105), .O(n11886));
  OAI112BHD U14813 ( .C1(n11879), .C2(_i_CLEFIA128_keyL _105), .A1(n11878), .B1(n8589), .O(n11884) );
  OA12EHD U14814 ( .B1(n11881), .B2(n11880), .A1(_i_CLEFIA128_state_reg _1), .O(n11883) );
  ND3EHD U14815 ( .I1(n11884), .I2(n11883), .I3(n11882), .O(n11885) );
  ND2DHD U14816 ( .I1(_i_CLEFIA128_keyK _45), .I2(_i_CLEFIA128_keyL _45), .O(n11888) );
  XOR2EHD U14817 ( .I1(_i_CLEFIA128_CON_T_xi _11), .I2(DOUT_109), .O(n11890));
  NR2CHD U14818 ( .I1(n12982), .I2(n12240), .O(n11909) );
  AN2EHD U14819 ( .I1(n9589), .I2(n6770), .O(n11912) );
  INVDHD U14820 ( .I(_i_CLEFIA128_keyK _46), .O(n14026) );
  INVDHD U14821 ( .I(_i_CLEFIA128_keyK _47), .O(n15353) );
  NR2CHD U14822 ( .I1(n15353), .I2(n14707), .O(n11924) );
  AN3EHD U14823 ( .I1(n8320), .I2(n9693), .I3(n13440), .O(n11933) );
  NR2CHD U14824 ( .I1(n13388), .I2(n12353), .O(n11940) );
  NR3BHD U14825 ( .I1(n11947), .I2(n13029), .I3(n13015), .O(n11953) );
  XOR2EHD U14826 ( .I1(_i_CLEFIA128_CON_T_x _3), .I2(DOUT_99), .O(n11969) );
  XNR2EHD U14827 ( .I1(_i_CLEFIA128_CON_T_reg_4 ), .I2(DOUT_101), .O(n11975));
  ND2KHD U14828 ( .I1(n12029), .I2(n12914), .O(n11991) );
  ND2DHD U14829 ( .I1(_i_CLEFIA128_keyK _34), .I2(_i_CLEFIA128_keyL _34), .O(n11984) );
  ND2DHD U14830 ( .I1(n8797), .I2(_i_CLEFIA128_keyK _34), .O(n11982) );
  OR3EHD U14831 ( .I1(n12006), .I2(n12005), .I3(n13605), .O(n12025) );
  INVDHD U14832 ( .I(_i_CLEFIA128_keyK _38), .O(n13802) );
  MXL2CHD U14833 ( .A(n12020), .B(n12019), .S(_i_CLEFIA128_keyL _38), .OB(n12021) );
  ND3CHD U14834 ( .I1(n12022), .I2(n12021), .I3(_i_CLEFIA128_state_reg _1), .O(n12023) );
  XNR2EHD U14835 ( .I1(n12024), .I2(n12023), .O(n12062) );
  ND2DHD U14836 ( .I1(n12915), .I2(n12031), .O(n12032) );
  NR2CHD U14837 ( .I1(n12260), .I2(n13150), .O(n12041) );
  ND2DHD U14838 ( .I1(n9603), .I2(n13602), .O(n12039) );
  INVDHD U14839 ( .I(n12062), .O(n12053) );
  ND2DHD U14840 ( .I1(n12030), .I2(n12044), .O(n12045) );
  NR3BHD U14841 ( .I1(n12047), .I2(n12046), .I3(n12277), .O(n12051) );
  NR2CHD U14842 ( .I1(n7550), .I2(n12049), .O(n12050) );
  ND2DHD U14843 ( .I1(n10095), .I2(n12901), .O(n12267) );
  ND2DHD U14844 ( .I1(n13121), .I2(n13130), .O(n12060) );
  ND2DHD U14845 ( .I1(n9807), .I2(n12171), .O(n12154) );
  ND3CHD U14846 ( .I1(n13512), .I2(n12296), .I3(n12154), .O(n12067) );
  ND2DHD U14847 ( .I1(n12298), .I2(n13510), .O(n13839) );
  OR3EHD U14848 ( .I1(n12068), .I2(n13839), .I3(n12067), .O(n12073) );
  OA13EHD U14849 ( .B1(n12074), .B2(n12073), .B3(n12072), .A1(n8294), .O(n12085) );
  INVDHD U14850 ( .I(n13682), .O(n12079) );
  ND2DHD U14851 ( .I1(n13646), .I2(n13838), .O(n13532) );
  INVDHD U14852 ( .I(n12075), .O(n12076) );
  ND2DHD U14853 ( .I1(n12145), .I2(n12076), .O(n13820) );
  ND3CHD U14854 ( .I1(n9098), .I2(n12306), .I3(n13820), .O(n12077) );
  NR2CHD U14855 ( .I1(n13532), .I2(n12077), .O(n12078) );
  ND3CHD U14856 ( .I1(n12079), .I2(n13814), .I3(n12078), .O(n12083) );
  AN2EHD U14857 ( .I1(n13810), .I2(n9741), .O(n12093) );
  INVDHD U14858 ( .I(n7165), .O(n12111) );
  NR2GHD U14859 ( .I1(n12111), .I2(n12898), .O(n12948) );
  AN2EHD U14860 ( .I1(n13592), .I2(n13589), .O(n12284) );
  INVDHD U14861 ( .I(n12905), .O(n12119) );
  NR2CHD U14862 ( .I1(n9674), .I2(n12120), .O(n12121) );
  AN2EHD U14863 ( .I1(n12128), .I2(n13130), .O(n12132) );
  NR2CHD U14864 ( .I1(n12129), .I2(n12902), .O(n12130) );
  INVDHD U14865 ( .I(n12133), .O(n12134) );
  AOI22BHD U14866 ( .A1(n15492), .A2(DIN_107), .B1(n7017), .B2(KEY_107), .O(n12142) );
  AN3EHD U14867 ( .I1(n6685), .I2(n12306), .I3(n12154), .O(n12157) );
  ND3CHD U14868 ( .I1(n12159), .I2(n9621), .I3(n13810), .O(n12160) );
  ND2DHD U14869 ( .I1(n13653), .I2(n13506), .O(n12169) );
  ND2DHD U14870 ( .I1(n7035), .I2(n12171), .O(n12174) );
  ND2DHD U14871 ( .I1(n8209), .I2(n7538), .O(n13537) );
  ND3CHD U14872 ( .I1(n12174), .I2(n13537), .I3(n13538), .O(n12175) );
  ND2DHD U14873 ( .I1(n12177), .I2(n12176), .O(n12178) );
  INVDHD U14874 ( .I(n13488), .O(n12180) );
  ND3CHD U14875 ( .I1(n12180), .I2(n13106), .I3(n13491), .O(n12184) );
  NR3BHD U14876 ( .I1(n12194), .I2(n13097), .I3(n12193), .O(n12197) );
  ND3CHD U14877 ( .I1(n12200), .I2(n12199), .I3(n12198), .O(n12201) );
  AN2EHD U14878 ( .I1(n8422), .I2(n13220), .O(n12204) );
  INVDHD U14879 ( .I(n12205), .O(n12206) );
  ND3CHD U14880 ( .I1(n12207), .I2(n12206), .I3(n13482), .O(n12213) );
  ND2DHD U14881 ( .I1(n8296), .I2(n12226), .O(n12219) );
  INVDHD U14882 ( .I(n12229), .O(n12230) );
  ND2HHD U14883 ( .I1(n12230), .I2(n13367), .O(n12231) );
  INVDHD U14884 ( .I(n12411), .O(n12239) );
  ND2DHD U14885 ( .I1(n13406), .I2(n9548), .O(n12242) );
  ND3CHD U14886 ( .I1(n12248), .I2(n9632), .I3(n13440), .O(n12250) );
  OAI12CHD U14887 ( .B1(n7830), .B2(n12251), .A1(n9676), .O(n12252) );
  ND2DHD U14888 ( .I1(n12902), .I2(n8228), .O(n12266) );
  AN3EHD U14889 ( .I1(n6543), .I2(n12267), .I3(n12266), .O(n12270) );
  AN2EHD U14890 ( .I1(n12268), .I2(n9772), .O(n12269) );
  INVDHD U14891 ( .I(n12272), .O(n12273) );
  ND2DHD U14892 ( .I1(n9772), .I2(n12276), .O(n13619) );
  NR3BHD U14893 ( .I1(n12279), .I2(n13172), .I3(n12395), .O(n12285) );
  NR2CHD U14894 ( .I1(n12282), .I2(n12281), .O(n12283) );
  ND2DHD U14895 ( .I1(n13005), .I2(n12335), .O(n12337) );
  ND2DHD U14896 ( .I1(n13448), .I2(n13004), .O(n12336) );
  ND3EHD U14897 ( .I1(n12343), .I2(n8320), .I3(n12369), .O(n12344) );
  ND2DHD U14898 ( .I1(n7830), .I2(n8296), .O(n12347) );
  ND2DHD U14899 ( .I1(n12414), .I2(n8394), .O(n12356) );
  ND2DHD U14900 ( .I1(n6930), .I2(n9676), .O(n13382) );
  ND2DHD U14901 ( .I1(n13448), .I2(n13382), .O(n12365) );
  OR3EHD U14902 ( .I1(n13446), .I2(n12365), .I3(n12967), .O(n12371) );
  INVDHD U14903 ( .I(n12374), .O(n12381) );
  INVDHD U14904 ( .I(n12377), .O(n13185) );
  ND2DHD U14905 ( .I1(n13185), .I2(n12915), .O(n13612) );
  ND3CHD U14906 ( .I1(n13121), .I2(n12917), .I3(n13612), .O(n12378) );
  ND2DHD U14907 ( .I1(n8185), .I2(n8228), .O(n12390) );
  ND2DHD U14908 ( .I1(n13128), .I2(n13627), .O(n12918) );
  OA13EHD U14909 ( .B1(n12397), .B2(n13140), .B3(n13631), .A1(n13634), .O(n12409) );
  ND2DHD U14910 ( .I1(n12402), .I2(n13614), .O(n12403) );
  OR2B1CHD U14911 ( .I1(n12411), .B1(n12410), .O(n12412) );
  ND2DHD U14912 ( .I1(n13448), .I2(n9679), .O(n12417) );
  ND2DHD U14913 ( .I1(n12424), .I2(n7037), .O(n13035) );
  AN3EHD U14914 ( .I1(n8433), .I2(n13000), .I3(n13019), .O(n12433) );
  AN2EHD U14915 ( .I1(n13036), .I2(n12436), .O(n12437) );
  AOI22BHD U14916 ( .A1(n15492), .A2(DIN_60), .B1(n7017), .B2(KEY_60), .O(n12446) );
  INVDHD U14917 ( .I(n12457), .O(n12458) );
  ND3CHD U14918 ( .I1(n12458), .I2(n8782), .I3(n12502), .O(n12459) );
  ND2DHD U14919 ( .I1(n12469), .I2(n12468), .O(n12471) );
  NR2CHD U14920 ( .I1(n12470), .I2(n12471), .O(n12472) );
  ND2DHD U14921 ( .I1(n6588), .I2(n12478), .O(n12482) );
  ND2DHD U14922 ( .I1(n8781), .I2(n9047), .O(n12481) );
  NR2CHD U14923 ( .I1(n12482), .I2(n12481), .O(n12490) );
  ND2DHD U14924 ( .I1(n12486), .I2(n12485), .O(n12488) );
  OR3EHD U14925 ( .I1(n12496), .I2(n12494), .I3(n12495), .O(n12509) );
  ND2DHD U14926 ( .I1(n12546), .I2(n12513), .O(n12514) );
  OAI112BHD U14927 ( .C1(n6839), .C2(n7128), .A1(n12519), .B1(n12623), .O(n12524) );
  INVDHD U14928 ( .I(n12633), .O(n12533) );
  OAI12CHD U14929 ( .B1(n12536), .B2(n12535), .A1(n12605), .O(n12550) );
  AN4CHD U14930 ( .I1(n9709), .I2(n12538), .I3(n12652), .I4(n12537), .O(n12543) );
  NR2CHD U14931 ( .I1(n12628), .I2(n12539), .O(n12542) );
  INVDHD U14932 ( .I(n12540), .O(n12541) );
  AN2EHD U14933 ( .I1(n9104), .I2(n12577), .O(n12554) );
  NR2CHD U14934 ( .I1(n12568), .I2(n12567), .O(n12569) );
  INVDHD U14935 ( .I(n12579), .O(n12580) );
  ND2DHD U14936 ( .I1(n9666), .I2(n12581), .O(n12584) );
  NR2CHD U14937 ( .I1(n12584), .I2(n12583), .O(n12589) );
  AOI22BHD U14938 ( .A1(n7045), .A2(n12595), .B1(n15504), .B2(n12594), .O(n12817) );
  AOI22BHD U14939 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _83), .B1(n15504), .B2(_i_CLEFIA128_keyK _19), .O(n12816) );
  INVDHD U14940 ( .I(n12596), .O(n12597) );
  NR2CHD U14941 ( .I1(n12599), .I2(n12600), .O(n12601) );
  INVDHD U14942 ( .I(n12620), .O(n12624) );
  INVDHD U14943 ( .I(n12626), .O(n12630) );
  NR2CHD U14944 ( .I1(n12628), .I2(n12627), .O(n12629) );
  NR2CHD U14945 ( .I1(n12634), .I2(n12633), .O(n12645) );
  NR2CHD U14946 ( .I1(n12636), .I2(n7138), .O(n12644) );
  ND2DHD U14947 ( .I1(n7154), .I2(n12637), .O(n12642) );
  ND3CHD U14948 ( .I1(n9663), .I2(n12640), .I3(n12639), .O(n12641) );
  INVDHD U14949 ( .I(n12650), .O(n12664) );
  NR2CHD U14950 ( .I1(n12654), .I2(n12653), .O(n12661) );
  AN3EHD U14951 ( .I1(n9663), .I2(n7154), .I3(n12657), .O(n12660) );
  INVDHD U14952 ( .I(n12658), .O(n12659) );
  ND3CHD U14953 ( .I1(n12660), .I2(n12661), .I3(n12659), .O(n12663) );
  ND2DHD U14954 ( .I1(n12669), .I2(n12668), .O(n12781) );
  ND3CHD U14955 ( .I1(n12678), .I2(n8564), .I3(n12708), .O(n12679) );
  AN2EHD U14956 ( .I1(n12869), .I2(n12689), .O(n12682) );
  NR2CHD U14957 ( .I1(n12684), .I2(n12683), .O(n12686) );
  ND2DHD U14958 ( .I1(n12690), .I2(n12689), .O(n12691) );
  INVDHD U14959 ( .I(n6970), .O(n12694) );
  AN3EHD U14960 ( .I1(n6706), .I2(n12714), .I3(n9735), .O(n12715) );
  XOR2EHD U14961 ( .I1(n12717), .I2(n12856), .O(n12718) );
  NR2CHD U14962 ( .I1(n12739), .I2(n12738), .O(n12741) );
  ND2DHD U14963 ( .I1(n12751), .I2(n9801), .O(n12753) );
  ND3CHD U14964 ( .I1(n12767), .I2(n12766), .I3(n12765), .O(n12774) );
  NR2CHD U14965 ( .I1(n12774), .I2(n12773), .O(n12775) );
  NR2CHD U14966 ( .I1(n12781), .I2(n12780), .O(n12782) );
  ND3CHD U14967 ( .I1(n12783), .I2(n12784), .I3(n8415), .O(n12785) );
  ND3CHD U14968 ( .I1(n12798), .I2(n12797), .I3(n8193), .O(n12803) );
  ND2DHD U14969 ( .I1(n12876), .I2(n8236), .O(n12801) );
  NR2EHD U14970 ( .I1(n12874), .I2(n12807), .O(n12812) );
  AOI22BHD U14971 ( .A1(n7017), .A2(KEY_19), .B1(n13292), .B2(n12818), .O(n12819) );
  OAI112BHD U14972 ( .C1(n10912), .C2(n12821), .A1(n12820), .B1(n12819), .O(n12823) );
  OAI22CHD U14973 ( .A1(n15488), .A2(n15513), .B1(n15512), .B2(n15491), .O(n12822) );
  ND2HHD U14974 ( .I1(n12825), .I2(n12824), .O(n6108) );
  ND2DHD U14975 ( .I1(n12830), .I2(n12829), .O(n12831) );
  ND3CHD U14976 ( .I1(n12833), .I2(n12832), .I3(n12831), .O(n12834) );
  OR2B1CHD U14977 ( .I1(n12836), .B1(n9723), .O(n12837) );
  NR2CHD U14978 ( .I1(n12839), .I2(n12838), .O(n12841) );
  ND2DHD U14979 ( .I1(n7155), .I2(n9723), .O(n12844) );
  NR2CHD U14980 ( .I1(n12849), .I2(n12848), .O(n12850) );
  NR2CHD U14981 ( .I1(n12852), .I2(n12851), .O(n12853) );
  AN2EHD U14982 ( .I1(n12878), .I2(n12856), .O(n12859) );
  ND3CHD U14983 ( .I1(n12859), .I2(n12858), .I3(n12857), .O(n12861) );
  NR2CHD U14984 ( .I1(n12861), .I2(n12860), .O(n12862) );
  ND2DHD U14985 ( .I1(n12866), .I2(n6670), .O(n12871) );
  ND2DHD U14986 ( .I1(n7155), .I2(n12868), .O(n12870) );
  NR2CHD U14987 ( .I1(n12871), .I2(n12870), .O(n12873) );
  ND2DHD U14988 ( .I1(n12873), .I2(n12872), .O(n12884) );
  AN3EHD U14989 ( .I1(n12877), .I2(n12878), .I3(n12876), .O(n12879) );
  ND3CHD U14990 ( .I1(n10207), .I2(n12879), .I3(n9590), .O(n12881) );
  AOI22BHD U14991 ( .A1(n7017), .A2(KEY_12), .B1(n13292), .B2(n12888), .O(n12889) );
  OAI112BHD U14992 ( .C1(n10912), .C2(n12891), .A1(n12890), .B1(n12889), .O(n12893) );
  OAI22CHD U14993 ( .A1(n15345), .A2(n15513), .B1(n15512), .B2(n15015), .O(n12892) );
  AOI22BHD U14994 ( .A1(n15492), .A2(DIN_124), .B1(n7017), .B2(KEY_124), .O(n12896) );
  OA12EHD U14995 ( .B1(n15499), .B2(n14321), .A1(n12896), .O(n12897) );
  ND3EHD U14996 ( .I1(n12899), .I2(n8175), .I3(n10294), .O(n13170) );
  ND2DHD U14997 ( .I1(n12900), .I2(n12901), .O(n12904) );
  ND2DHD U14998 ( .I1(n12902), .I2(n8223), .O(n12903) );
  ND3CHD U14999 ( .I1(n13183), .I2(n12904), .I3(n12903), .O(n12907) );
  ND2DHD U15000 ( .I1(n12905), .I2(n9639), .O(n12906) );
  ND3CHD U15001 ( .I1(n12908), .I2(n12909), .I3(n12910), .O(n12911) );
  ND3CHD U15002 ( .I1(n12915), .I2(n8897), .I3(n9777), .O(n12916) );
  ND2DHD U15003 ( .I1(n13194), .I2(n12916), .O(n12919) );
  ND3CHD U15004 ( .I1(n12925), .I2(n12924), .I3(n12923), .O(n12926) );
  ND2DHD U15005 ( .I1(n12928), .I2(n12929), .O(n12940) );
  ND3CHD U15006 ( .I1(n12933), .I2(n9463), .I3(n12934), .O(n12938) );
  AN2EHD U15007 ( .I1(n13187), .I2(n12945), .O(n12946) );
  AN3EHD U15008 ( .I1(n12946), .I2(n13182), .I3(n7031), .O(n12947) );
  ND2DHD U15009 ( .I1(n12950), .I2(n13427), .O(n12954) );
  ND2DHD U15010 ( .I1(n8784), .I2(n7830), .O(n12963) );
  INVDHD U15011 ( .I(n12981), .O(n12994) );
  INVDHD U15012 ( .I(n12982), .O(n12987) );
  ND2DHD U15013 ( .I1(n8214), .I2(n8229), .O(n12983) );
  NR2CHD U15014 ( .I1(n12985), .I2(n12984), .O(n12986) );
  ND3CHD U15015 ( .I1(n6980), .I2(n13001), .I3(n13000), .O(n13003) );
  ND3CHD U15016 ( .I1(n13019), .I2(n13018), .I3(n13371), .O(n13020) );
  AN2EHD U15017 ( .I1(n13022), .I2(n13021), .O(n13023) );
  ND3CHD U15018 ( .I1(n13023), .I2(n9093), .I3(n13024), .O(n13027) );
  NR2CHD U15019 ( .I1(n13034), .I2(n13033), .O(n13038) );
  AN3EHD U15020 ( .I1(n9084), .I2(n13036), .I3(n13035), .O(n13037) );
  XNR2KHD U15021 ( .I1(n14367), .I2(n13040), .O(n15134) );
  AOI22BHD U15022 ( .A1(n7017), .A2(KEY_82), .B1(n13292), .B2(n13042), .O(n13043) );
  OAI112BHD U15023 ( .C1(n10912), .C2(n13045), .A1(n13044), .B1(n13043), .O(n13047) );
  OAI22CHD U15024 ( .A1(n14904), .A2(n15513), .B1(n15512), .B2(n15130), .O(n13046) );
  AN2HHD U15025 ( .I1(n13051), .I2(n13050), .O(n13052) );
  ND2DHD U15026 ( .I1(n14081), .I2(n13479), .O(n13059) );
  ND3CHD U15027 ( .I1(n9605), .I2(n13478), .I3(n13085), .O(n13086) );
  NR2CHD U15028 ( .I1(n13086), .I2(n13087), .O(n13093) );
  NR2CHD U15029 ( .I1(n13090), .I2(n13089), .O(n13091) );
  ND2DHD U15030 ( .I1(n9184), .I2(n13100), .O(n13101) );
  OAI12CHD U15031 ( .B1(n13109), .B2(n13108), .A1(n9537), .O(n13113) );
  ND2DHD U15032 ( .I1(n13132), .I2(n8228), .O(n13133) );
  AN3EHD U15033 ( .I1(n13142), .I2(n13182), .I3(n13614), .O(n13148) );
  INVDHD U15034 ( .I(n13152), .O(n13154) );
  ND3CHD U15035 ( .I1(n13153), .I2(n13155), .I3(n13154), .O(n13156) );
  AOI22BHD U15036 ( .A1(n15492), .A2(DIN_122), .B1(n7017), .B2(KEY_122), .O(n13162) );
  OAI12CHD U15037 ( .B1(n15499), .B2(n15337), .A1(n13162), .O(n13163) );
  NR2CHD U15038 ( .I1(n13166), .I2(n13165), .O(n13167) );
  NR2CHD U15039 ( .I1(n13174), .I2(n13173), .O(n13180) );
  INVDHD U15040 ( .I(n13175), .O(n13177) );
  NR2CHD U15041 ( .I1(n13177), .I2(n13176), .O(n13178) );
  ND2DHD U15042 ( .I1(n12030), .I2(n13185), .O(n13186) );
  ND3CHD U15043 ( .I1(n13188), .I2(n13187), .I3(n13186), .O(n13189) );
  NR2GHD U15044 ( .I1(n13189), .I2(n13190), .O(n13621) );
  ND2DHD U15045 ( .I1(n8183), .I2(n8223), .O(n13198) );
  INVDHD U15046 ( .I(n13576), .O(n13200) );
  ND2DHD U15047 ( .I1(n13204), .I2(n13203), .O(n13205) );
  ND2DHD U15048 ( .I1(n9886), .I2(n13207), .O(n13210) );
  ND2DHD U15049 ( .I1(n13223), .I2(n13222), .O(n13225) );
  NR2CHD U15050 ( .I1(n13227), .I2(n13226), .O(n13228) );
  ND2DHD U15051 ( .I1(n6932), .I2(n13246), .O(n13248) );
  NR2CHD U15052 ( .I1(n13248), .I2(n13247), .O(n13249) );
  AOI22BHD U15053 ( .A1(n7017), .A2(KEY_68), .B1(n13292), .B2(n13257), .O(n13258) );
  OAI112BHD U15054 ( .C1(n10912), .C2(n13260), .A1(n13259), .B1(n13258), .O(n13262) );
  OAI22CHD U15055 ( .A1(n14983), .A2(n15513), .B1(n15512), .B2(n14814), .O(n13261) );
  OAI112BHD U15056 ( .C1(n14837), .C2(n13265), .A1(n13264), .B1(n13263), .O(n6154) );
  OAI112BHD U15057 ( .C1(n13272), .C2(n10912), .A1(n13271), .B1(n13270), .O(n13273) );
  AOI12CHD U15058 ( .B1(n10928), .B2(DOUT_3), .A1(n13273), .O(n13275) );
  ND2HHD U15059 ( .I1(n14721), .I2(n13284), .O(n13285) );
  BUFQHD U15060 ( .I(n13285), .O(n15416) );
  ND2DHD U15061 ( .I1(n13291), .I2(n13287), .O(n13288) );
  ND3EHD U15062 ( .I1(n15420), .I2(n15416), .I3(n13293), .O(n14796) );
  OAI112BHD U15063 ( .C1(n13277), .C2(n14934), .A1(n13295), .B1(n13294), .O(n6232) );
  OAI112BHD U15064 ( .C1(n13277), .C2(n15212), .A1(n13299), .B1(n13298), .O(n6242) );
  OAI112BHD U15065 ( .C1(n13277), .C2(n15300), .A1(n13303), .B1(n13302), .O(n6233) );
  OAI112BHD U15066 ( .C1(n13277), .C2(n15263), .A1(n13307), .B1(n13306), .O(n6245) );
  OAI112BHD U15067 ( .C1(n13277), .C2(n14991), .A1(n13311), .B1(n13310), .O(n6240) );
  OAI112BHD U15068 ( .C1(n13277), .C2(n15209), .A1(n13315), .B1(n13314), .O(n6235) );
  OAI112BHD U15069 ( .C1(n13277), .C2(n8902), .A1(n13319), .B1(n13318), .O(n6298) );
  OAI112BHD U15070 ( .C1(n13277), .C2(n15069), .A1(n13323), .B1(n13322), .O(n6297) );
  OAI112BHD U15071 ( .C1(n13277), .C2(n9528), .A1(n13327), .B1(n13326), .O(n6291) );
  OAI112BHD U15072 ( .C1(n13277), .C2(n15304), .A1(n13331), .B1(n13330), .O(n6226) );
  OAI112BHD U15073 ( .C1(n13277), .C2(n14988), .A1(n13335), .B1(n13334), .O(n6247) );
  OAI112BHD U15074 ( .C1(n13277), .C2(n15064), .A1(n13338), .B1(n8386), .O(n6224) );
  OAI112BHD U15075 ( .C1(n13277), .C2(n15089), .A1(n13343), .B1(n13342), .O(n6294) );
  OAI112BHD U15076 ( .C1(n13277), .C2(n14931), .A1(n13347), .B1(n13346), .O(n6225) );
  OAI112BHD U15077 ( .C1(n13277), .C2(n15189), .A1(n13351), .B1(n13350), .O(n6292) );
  OAI112BHD U15078 ( .C1(n13277), .C2(n15408), .A1(n13359), .B1(n13358), .O(n6229) );
  XNR2EHD U15079 ( .I1(DOUT_22), .I2(n14489), .O(n13360) );
  AOI22BHD U15080 ( .A1(n15492), .A2(DIN_118), .B1(n7017), .B2(KEY_118), .O(n13361) );
  INVDHD U15081 ( .I(n13444), .O(n13362) );
  ND3CHD U15082 ( .I1(n13366), .I2(n13365), .I3(n9084), .O(n13368) );
  ND2DHD U15083 ( .I1(n13370), .I2(n13369), .O(n13378) );
  ND3CHD U15084 ( .I1(n13373), .I2(n13372), .I3(n13371), .O(n13374) );
  OR2B1CHD U15085 ( .I1(n13376), .B1(n13428), .O(n13377) );
  ND2DHD U15086 ( .I1(n9632), .I2(n13382), .O(n13385) );
  ND2DHD U15087 ( .I1(n6770), .I2(n9548), .O(n13384) );
  ND2DHD U15088 ( .I1(n13387), .I2(n13386), .O(n13393) );
  AN3EHD U15089 ( .I1(n13394), .I2(n13409), .I3(n13395), .O(n13415) );
  ND2DHD U15090 ( .I1(n13457), .I2(n13397), .O(n13403) );
  ND3CHD U15091 ( .I1(n13400), .I2(n13402), .I3(n9589), .O(n13466) );
  NR2CHD U15092 ( .I1(n13403), .I2(n13466), .O(n13405) );
  ND2DHD U15093 ( .I1(n13404), .I2(n13405), .O(n13412) );
  NR2CHD U15094 ( .I1(n13407), .I2(n13408), .O(n13410) );
  ND2DHD U15095 ( .I1(n13410), .I2(n13409), .O(n13411) );
  OA22EHD U15096 ( .A1(n13415), .A2(n13416), .B1(n13414), .B2(n13413), .O(n13417) );
  NR2CHD U15097 ( .I1(n13423), .I2(n13422), .O(n13424) );
  ND2DHD U15098 ( .I1(n13448), .I2(n13447), .O(n13450) );
  NR2CHD U15099 ( .I1(n13449), .I2(n13450), .O(n13451) );
  ND3CHD U15100 ( .I1(n13457), .I2(n9574), .I3(n9093), .O(n13465) );
  XNR2EHD U15101 ( .I1(DOUT_86), .I2(n9664), .O(n13501) );
  INVDHD U15102 ( .I(n13477), .O(n13486) );
  ND3CHD U15103 ( .I1(n13479), .I2(n13478), .I3(n7077), .O(n13481) );
  ND3CHD U15104 ( .I1(n13483), .I2(n13482), .I3(n14065), .O(n13484) );
  ND2DHD U15105 ( .I1(n8250), .I2(n8197), .O(n13496) );
  OAI13BHD U15106 ( .B1(n13497), .B2(n13498), .B3(n10297), .A1(n14067), .O(n13499) );
  XOR2HHD U15107 ( .I1(n9370), .I2(n14106), .O(n13500) );
  ND2DHD U15108 ( .I1(n15178), .I2(n15500), .O(n13502) );
  ND3CHD U15109 ( .I1(n13504), .I2(n13503), .I3(n13502), .O(n6212) );
  XNR3EHD U15110 ( .I1(DOUT_25), .I2(n6889), .I3(n7789), .O(n13505) );
  XNR2EHD U15111 ( .I1(n14144), .I2(n13505), .O(n15468) );
  NR2CHD U15112 ( .I1(n13654), .I2(n13507), .O(n13508) );
  ND2DHD U15113 ( .I1(n13509), .I2(n13508), .O(n13520) );
  ND2DHD U15114 ( .I1(n13513), .I2(n13512), .O(n13515) );
  ND2DHD U15115 ( .I1(n13516), .I2(n13533), .O(n13517) );
  OR3EHD U15116 ( .I1(n13682), .I2(n13518), .I3(n13517), .O(n13519) );
  ND2DHD U15117 ( .I1(n6872), .I2(n8279), .O(n13522) );
  OR3EHD U15118 ( .I1(n13682), .I2(n13540), .I3(n13679), .O(n13545) );
  ND2DHD U15119 ( .I1(n13642), .I2(n13541), .O(n13542) );
  NR2CHD U15120 ( .I1(n13542), .I2(n9299), .O(n13543) );
  ND2DHD U15121 ( .I1(n13823), .I2(n13543), .O(n13544) );
  AN2EHD U15122 ( .I1(n13659), .I2(n13810), .O(n13546) );
  ND3CHD U15123 ( .I1(n13546), .I2(n13838), .I3(n6582), .O(n13548) );
  OR3EHD U15124 ( .I1(n13549), .I2(n13548), .I3(n13547), .O(n13552) );
  XNR3EHD U15125 ( .I1(DOUT_89), .I2(n8870), .I3(n9705), .O(n13557) );
  ND2DHD U15126 ( .I1(n14913), .I2(n15500), .O(n13560) );
  AOI22BHD U15127 ( .A1(n15492), .A2(DIN_121), .B1(n7017), .B2(KEY_121), .O(n13558) );
  ND3CHD U15128 ( .I1(n13561), .I2(n13560), .I3(n13559), .O(n6215) );
  AOI22BHD U15129 ( .A1(n15492), .A2(DIN_57), .B1(n7017), .B2(KEY_57), .O(n13562) );
  ND3CHD U15130 ( .I1(n13565), .I2(n13564), .I3(n13563), .O(n6183) );
  ND2DHD U15131 ( .I1(n14813), .I2(n15500), .O(n13569) );
  AOI22BHD U15132 ( .A1(n15492), .A2(DIN_54), .B1(n7017), .B2(KEY_54), .O(n13566) );
  ND3CHD U15133 ( .I1(n13569), .I2(n13568), .I3(n13567), .O(n6180) );
  AOI22BHD U15134 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _126), .B1(n15504), .B2(_i_CLEFIA128_keyK _62), .O(n13691) );
  NR3BHD U15135 ( .I1(n13576), .I2(n13574), .I3(n13575), .O(n13581) );
  NR2CHD U15136 ( .I1(n13579), .I2(n13578), .O(n13580) );
  INVDHD U15137 ( .I(n13582), .O(n13583) );
  ND2DHD U15138 ( .I1(n13590), .I2(n13589), .O(n13599) );
  ND2DHD U15139 ( .I1(n13592), .I2(n9603), .O(n13598) );
  ND3CHD U15140 ( .I1(n13596), .I2(n13595), .I3(n13594), .O(n13597) );
  NR3BHD U15141 ( .I1(n13599), .I2(n13598), .I3(n13597), .O(n13600) );
  ND3CHD U15142 ( .I1(n13607), .I2(n8410), .I3(n13606), .O(n13609) );
  OR3EHD U15143 ( .I1(n13616), .I2(n13617), .I3(n13615), .O(n13625) );
  OA13EHD U15144 ( .B1(n13623), .B2(n13624), .B3(n13625), .A1(n13622), .O(n13639) );
  INVDHD U15145 ( .I(n13626), .O(n13633) );
  AN3EHD U15146 ( .I1(n9886), .I2(n6543), .I3(n13627), .O(n13630) );
  OA13EHD U15147 ( .B1(n13637), .B2(n9878), .B3(n13635), .A1(n13634), .O(n13638) );
  NR2CHD U15148 ( .I1(n13648), .I2(n13647), .O(n13649) );
  ND3CHD U15149 ( .I1(n13660), .I2(n13659), .I3(n9094), .O(n13665) );
  OR2B1CHD U15150 ( .I1(n13662), .B1(n13661), .O(n13664) );
  OA13EHD U15151 ( .B1(n13666), .B2(n13667), .B3(n13816), .A1(n13826), .O(n13668) );
  AN2B1CHD U15152 ( .I1(n9098), .B1(n13670), .O(n13672) );
  ND2DHD U15153 ( .I1(n13673), .I2(n13823), .O(n13674) );
  ND3CHD U15154 ( .I1(n13677), .I2(n9814), .I3(n8758), .O(n13678) );
  ND3CHD U15155 ( .I1(n13685), .I2(n13684), .I3(n6684), .O(n13686) );
  OA13EHD U15156 ( .B1(n13687), .B2(n13686), .B3(n13848), .A1(n13817), .O(n13688) );
  AOI22BHD U15157 ( .A1(n7017), .A2(KEY_94), .B1(n13292), .B2(n13692), .O(n13693) );
  OAI112BHD U15158 ( .C1(n10912), .C2(n13695), .A1(n13694), .B1(n13693), .O(n13697) );
  OAI22CHD U15159 ( .A1(n15494), .A2(n15513), .B1(n15512), .B2(n15498), .O(n13696) );
  AOI22BHD U15160 ( .A1(n7045), .A2(n13700), .B1(n15504), .B2(n13699), .O(n13704) );
  AOI22BHD U15161 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _88), .B1(n15504), .B2(_i_CLEFIA128_keyK _24), .O(n13703) );
  XOR2EHD U15162 ( .I1(DOUT_24), .I2(n9657), .O(n13702) );
  AOI22BHD U15163 ( .A1(n7017), .A2(KEY_24), .B1(n13292), .B2(n13705), .O(n13706) );
  OAI112BHD U15164 ( .C1(n10912), .C2(n13708), .A1(n13707), .B1(n13706), .O(n13710) );
  OAI22CHD U15165 ( .A1(n14608), .A2(n15513), .B1(n15512), .B2(n14880), .O(n13709) );
  AOI22BHD U15166 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _65), .B1(n15504), .B2(_i_CLEFIA128_keyK _1), .O(n13719) );
  AOI22BHD U15167 ( .A1(n7045), .A2(n13714), .B1(n15504), .B2(n13713), .O(n13718) );
  MUX2EHD U15168 ( .A(n13719), .B(n13718), .S(n15200), .O(n13727) );
  AOI22BHD U15169 ( .A1(n7017), .A2(KEY_1), .B1(n13292), .B2(n13720), .O(n13721) );
  OAI112BHD U15170 ( .C1(n10912), .C2(n13723), .A1(n13722), .B1(n13721), .O(n13725) );
  OAI22CHD U15171 ( .A1(n15271), .A2(n15513), .B1(n15512), .B2(n15258), .O(n13724) );
  NR2CHD U15172 ( .I1(n13725), .I2(n13724), .O(n13726) );
  AOI22BHD U15173 ( .A1(n7045), .A2(n13729), .B1(n15504), .B2(n13728), .O(n13733) );
  AOI22BHD U15174 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _81), .B1(n15504), .B2(_i_CLEFIA128_keyK _17), .O(n13732) );
  XOR2EHD U15175 ( .I1(DOUT_17), .I2(n8309), .O(n13731) );
  AOI22BHD U15176 ( .A1(n7017), .A2(KEY_17), .B1(n13292), .B2(n13734), .O(n13735) );
  OAI112BHD U15177 ( .C1(n10912), .C2(n13737), .A1(n13736), .B1(n13735), .O(n13739) );
  OAI22CHD U15178 ( .A1(n14871), .A2(n15513), .B1(n15512), .B2(n15141), .O(n13738) );
  NR2CHD U15179 ( .I1(n13739), .I2(n13738), .O(n13740) );
  XNR3EHD U15180 ( .I1(DOUT_64), .I2(n9775), .I3(n14996), .O(n13743) );
  ND2DHD U15181 ( .I1(n15152), .I2(n15500), .O(n13746) );
  AOI22BHD U15182 ( .A1(n15492), .A2(DIN_96), .B1(n7017), .B2(KEY_96), .O(n13744) );
  ND3CHD U15183 ( .I1(n13747), .I2(n13746), .I3(n13745), .O(n6190) );
  ND2DHD U15184 ( .I1(n15520), .I2(n15500), .O(n13751) );
  ND2DHD U15185 ( .I1(n15152), .I2(n11130), .O(n13750) );
  AOI22BHD U15186 ( .A1(n15492), .A2(DIN_32), .B1(n7017), .B2(KEY_32), .O(n13748) );
  ND3CHD U15187 ( .I1(n13751), .I2(n13750), .I3(n13749), .O(n6221) );
  AOI22BHD U15188 ( .A1(n7045), .A2(n9974), .B1(n15504), .B2(n13752), .O(n13756) );
  AOI22BHD U15189 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _73), .B1(n15504), .B2(_i_CLEFIA128_keyK _9), .O(n13755) );
  AOI22BHD U15190 ( .A1(n7017), .A2(KEY_9), .B1(n13292), .B2(n13757), .O(n13758) );
  OAI112BHD U15191 ( .C1(n10912), .C2(n13760), .A1(n13759), .B1(n13758), .O(n13762) );
  OAI22CHD U15192 ( .A1(n15106), .A2(n15450), .B1(n15512), .B2(n15115), .O(n13761) );
  NR2CHD U15193 ( .I1(n13762), .I2(n13761), .O(n13763) );
  AOI22BHD U15194 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _119), .B1(n15504), .B2(_i_CLEFIA128_keyK _55), .O(n13769) );
  XNR2EHD U15195 ( .I1(DOUT_87), .I2(n8786), .O(n13768) );
  AOI22BHD U15196 ( .A1(n7017), .A2(KEY_87), .B1(n13292), .B2(n13770), .O(n13771) );
  OAI112BHD U15197 ( .C1(n10912), .C2(n13773), .A1(n13772), .B1(n13771), .O(n13775) );
  OAI22CHD U15198 ( .A1(n15432), .A2(n15450), .B1(n15512), .B2(n15437), .O(n13774) );
  AOI22BHD U15199 ( .A1(n7045), .A2(n13778), .B1(n15504), .B2(n13777), .O(n13781) );
  AOI22BHD U15200 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _80), .B1(n15504), .B2(_i_CLEFIA128_keyK _16), .O(n13780) );
  AOI22BHD U15201 ( .A1(n7017), .A2(KEY_16), .B1(n13292), .B2(n13782), .O(n13783) );
  OAI112BHD U15202 ( .C1(n10912), .C2(n13785), .A1(n13784), .B1(n13783), .O(n13787) );
  OAI22CHD U15203 ( .A1(n15369), .A2(n15450), .B1(n15512), .B2(n15373), .O(n13786) );
  NR2CHD U15204 ( .I1(n13787), .I2(n13786), .O(n13788) );
  AOI22BHD U15205 ( .A1(n7045), .A2(n13791), .B1(n15504), .B2(n13790), .O(n13793) );
  AOI22BHD U15206 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _95), .B1(n15504), .B2(_i_CLEFIA128_keyK _31), .O(n13792) );
  AOI22BHD U15207 ( .A1(n7017), .A2(KEY_31), .B1(n13292), .B2(n13794), .O(n13795) );
  OAI112BHD U15208 ( .C1(n10912), .C2(n13797), .A1(n13796), .B1(n13795), .O(n13799) );
  OAI22CHD U15209 ( .A1(n15417), .A2(n15513), .B1(n15512), .B2(n14866), .O(n13798) );
  NR2CHD U15210 ( .I1(n13799), .I2(n13798), .O(n13800) );
  AOI22BHD U15211 ( .A1(n7045), .A2(n13803), .B1(n15504), .B2(n13802), .O(n13853) );
  ND2DHD U15212 ( .I1(n13829), .I2(n9621), .O(n13831) );
  AN2B1CHD U15213 ( .I1(n13837), .B1(n13836), .O(n13847) );
  NR2CHD U15214 ( .I1(n13840), .I2(n13839), .O(n13846) );
  AN3EHD U15215 ( .I1(n13842), .I2(n13844), .I3(n13843), .O(n13845) );
  ND3CHD U15216 ( .I1(n13847), .I2(n13846), .I3(n13845), .O(n13849) );
  AOI22BHD U15217 ( .A1(n7017), .A2(KEY_70), .B1(n13292), .B2(n13854), .O(n13855) );
  OAI112BHD U15218 ( .C1(n10912), .C2(n13857), .A1(n13856), .B1(n13855), .O(n13859) );
  OAI22CHD U15219 ( .A1(n15442), .A2(n15450), .B1(n15512), .B2(n15428), .O(n13858) );
  NR2CHD U15220 ( .I1(n13859), .I2(n13858), .O(n13860) );
  ND2DHD U15221 ( .I1(n15392), .I2(n11130), .O(n13864) );
  AOI22BHD U15222 ( .A1(n15492), .A2(DIN_104), .B1(n7017), .B2(KEY_104), .O(n13861) );
  ND3CHD U15223 ( .I1(n13864), .I2(n13863), .I3(n13862), .O(n6198) );
  ND2DHD U15224 ( .I1(n15392), .I2(n15500), .O(n13868) );
  AOI22BHD U15225 ( .A1(n15492), .A2(DIN_40), .B1(n7017), .B2(KEY_40), .O(n13865) );
  OA12EHD U15226 ( .B1(n15499), .B2(n15385), .A1(n13865), .O(n13867) );
  ND2DHD U15227 ( .I1(n15193), .I2(n11130), .O(n13866) );
  AOI22BHD U15228 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _90), .B1(n15504), .B2(_i_CLEFIA128_keyK _26), .O(n13872) );
  AOI22BHD U15229 ( .A1(n7045), .A2(n13870), .B1(n15504), .B2(n13869), .O(n13871) );
  AOI22BHD U15230 ( .A1(n7017), .A2(KEY_26), .B1(n13292), .B2(n13873), .O(n13874) );
  OAI112BHD U15231 ( .C1(n10912), .C2(n13876), .A1(n13875), .B1(n13874), .O(n13878) );
  OAI22CHD U15232 ( .A1(n15337), .A2(n15513), .B1(n15512), .B2(n14959), .O(n13877) );
  AOI22BHD U15233 ( .A1(n7045), .A2(n13882), .B1(n15504), .B2(n13881), .O(n13885) );
  AOI22BHD U15234 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _87), .B1(n15504), .B2(_i_CLEFIA128_keyK _23), .O(n13884) );
  XNR2EHD U15235 ( .I1(n13911), .I2(n8774), .O(n13883) );
  AOI22BHD U15236 ( .A1(n7017), .A2(KEY_23), .B1(n13292), .B2(n13886), .O(n13887) );
  OAI112BHD U15237 ( .C1(n10912), .C2(n13889), .A1(n13888), .B1(n13887), .O(n13891) );
  OAI22CHD U15238 ( .A1(n15437), .A2(n15513), .B1(n15512), .B2(n15432), .O(n13890) );
  NR2CHD U15239 ( .I1(n13891), .I2(n13890), .O(n13892) );
  AOI22BHD U15240 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _82), .B1(n15504), .B2(_i_CLEFIA128_keyK _18), .O(n13900) );
  AOI22BHD U15241 ( .A1(n7045), .A2(n13894), .B1(n15504), .B2(n13893), .O(n13899) );
  XOR2HHD U15242 ( .I1(n13898), .I2(n13897), .O(n15131) );
  AOI22BHD U15243 ( .A1(n7017), .A2(KEY_18), .B1(n13292), .B2(n13901), .O(n13902) );
  OAI112BHD U15244 ( .C1(n10912), .C2(n13904), .A1(n13903), .B1(n13902), .O(n13906) );
  OAI22CHD U15245 ( .A1(n15130), .A2(n15513), .B1(n15512), .B2(n14904), .O(n13905) );
  NR2CHD U15246 ( .I1(n13906), .I2(n13905), .O(n13907) );
  AOI22BHD U15247 ( .A1(n7045), .A2(n13910), .B1(n15504), .B2(n13909), .O(n13914) );
  AOI22BHD U15248 ( .A1(n7017), .A2(KEY_30), .B1(n13292), .B2(n13915), .O(n13916) );
  OAI112BHD U15249 ( .C1(n10912), .C2(n13918), .A1(n13917), .B1(n13916), .O(n13920) );
  OAI22CHD U15250 ( .A1(n15498), .A2(n15513), .B1(n15512), .B2(n15494), .O(n13919) );
  NR2CHD U15251 ( .I1(n13920), .I2(n13919), .O(n13921) );
  AOI22BHD U15252 ( .A1(n7045), .A2(n7575), .B1(n15504), .B2(n13922), .O(n13928) );
  XNR3EHD U15253 ( .I1(n7789), .I2(n13924), .I3(n13923), .O(n13925) );
  AOI22BHD U15254 ( .A1(n7017), .A2(KEY_2), .B1(n13292), .B2(n13929), .O(n13930) );
  OAI112BHD U15255 ( .C1(n10912), .C2(n13932), .A1(n13931), .B1(n13930), .O(n13934) );
  OAI22CHD U15256 ( .A1(n15329), .A2(n15450), .B1(n15512), .B2(n15330), .O(n13933) );
  NR2CHD U15257 ( .I1(n13934), .I2(n13933), .O(n13935) );
  AOI22BHD U15258 ( .A1(n7045), .A2(n13937), .B1(n15504), .B2(n13936), .O(n13940) );
  AOI22BHD U15259 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _112), .B1(n15504), .B2(_i_CLEFIA128_keyK _48), .O(n13939) );
  XOR3EHD U15260 ( .I1(DOUT_80), .I2(n9775), .I3(n8870), .O(n13938) );
  AOI22BHD U15261 ( .A1(n7017), .A2(KEY_80), .B1(n13292), .B2(n13941), .O(n13942) );
  OAI112BHD U15262 ( .C1(n10912), .C2(n13944), .A1(n13943), .B1(n13942), .O(n13946) );
  OAI22CHD U15263 ( .A1(n15373), .A2(n15513), .B1(n15512), .B2(n15369), .O(n13945) );
  NR2CHD U15264 ( .I1(n13946), .I2(n13945), .O(n13947) );
  XOR2EHD U15265 ( .I1(DOUT_14), .I2(n9960), .O(n13953) );
  XOR2HHD U15266 ( .I1(n7256), .I2(n6808), .O(n13952) );
  AOI22BHD U15267 ( .A1(n7017), .A2(KEY_14), .B1(n13292), .B2(n13954), .O(n13955) );
  OAI112BHD U15268 ( .C1(n10912), .C2(n13957), .A1(n13956), .B1(n13955), .O(n13959) );
  OAI22CHD U15269 ( .A1(n15452), .A2(n15450), .B1(n15512), .B2(n15446), .O(n13958) );
  AOI22BHD U15270 ( .A1(n15492), .A2(DIN_111), .B1(n7017), .B2(KEY_111), .O(n13962) );
  XOR2EHD U15271 ( .I1(n9775), .I2(n7935), .O(n13964) );
  XOR2EHD U15272 ( .I1(DOUT_79), .I2(n9370), .O(n13963) );
  AOI22BHD U15273 ( .A1(n15492), .A2(DIN_47), .B1(n7017), .B2(KEY_47), .O(n13966) );
  AOI22BHD U15274 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _74), .B1(n15504), .B2(_i_CLEFIA128_keyK _10), .O(n13975) );
  AOI22BHD U15275 ( .A1(n7045), .A2(n13971), .B1(n15504), .B2(n13970), .O(n13974) );
  AOI22BHD U15276 ( .A1(n7017), .A2(KEY_10), .B1(n13292), .B2(n13976), .O(n13977) );
  OAI112BHD U15277 ( .C1(n10912), .C2(n13979), .A1(n13978), .B1(n13977), .O(n13981) );
  OAI22CHD U15278 ( .A1(n15393), .A2(n15513), .B1(n15512), .B2(n14802), .O(n13980) );
  AOI22BHD U15279 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _86), .B1(n15504), .B2(_i_CLEFIA128_keyK _22), .O(n13987) );
  AOI22BHD U15280 ( .A1(n7017), .A2(KEY_22), .B1(n13292), .B2(n13988), .O(n13989) );
  OAI112BHD U15281 ( .C1(n10912), .C2(n13991), .A1(n13990), .B1(n13989), .O(n13993) );
  OAI22CHD U15282 ( .A1(n15251), .A2(n15513), .B1(n15512), .B2(n15286), .O(n13992) );
  NR2CHD U15283 ( .I1(n13993), .I2(n13992), .O(n13994) );
  AOI22BHD U15284 ( .A1(n7017), .A2(KEY_86), .B1(n13292), .B2(n13997), .O(n13998) );
  OAI112BHD U15285 ( .C1(n10912), .C2(n14000), .A1(n13999), .B1(n13998), .O(n14002) );
  OAI22CHD U15286 ( .A1(n15286), .A2(n15450), .B1(n15512), .B2(n15251), .O(n14001) );
  AOI22BHD U15287 ( .A1(n15492), .A2(DIN_127), .B1(n7017), .B2(KEY_127), .O(n14004) );
  OAI12CHD U15288 ( .B1(n15499), .B2(n15417), .A1(n14004), .O(n14009) );
  NR2CHD U15289 ( .I1(n15512), .I2(n14525), .O(n14008) );
  OR3EHD U15290 ( .I1(n14009), .I2(n14008), .I3(n14007), .O(n6349) );
  AOI22BHD U15291 ( .A1(n15492), .A2(DIN_63), .B1(n7017), .B2(KEY_63), .O(n14010) );
  AOI22BHD U15292 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _70), .B1(n15504), .B2(_i_CLEFIA128_keyK _6), .O(n14018) );
  XOR2EHD U15293 ( .I1(DOUT_6), .I2(n8774), .O(n14017) );
  AOI22BHD U15294 ( .A1(n7017), .A2(KEY_6), .B1(n13292), .B2(n14019), .O(n14020) );
  OAI112BHD U15295 ( .C1(n10912), .C2(n14022), .A1(n14021), .B1(n14020), .O(n14024) );
  OAI22CHD U15296 ( .A1(n15428), .A2(n15450), .B1(n15512), .B2(n15442), .O(n14023) );
  AOI22BHD U15297 ( .A1(n7045), .A2(n14027), .B1(n15504), .B2(n14026), .O(n14032) );
  AOI22BHD U15298 ( .A1(n7017), .A2(KEY_78), .B1(n13292), .B2(n14033), .O(n14034) );
  OAI112BHD U15299 ( .C1(n10912), .C2(n14036), .A1(n14035), .B1(n14034), .O(n14038) );
  OAI22CHD U15300 ( .A1(n15446), .A2(n15513), .B1(n15512), .B2(n15452), .O(n14037) );
  AOI22BHD U15301 ( .A1(n7045), .A2(n14041), .B1(n15504), .B2(n14040), .O(n14093) );
  AOI22BHD U15302 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _120), .B1(n15504), .B2(_i_CLEFIA128_keyK _56), .O(n14092) );
  INVDHD U15303 ( .I(n14048), .O(n14050) );
  ND2DHD U15304 ( .I1(n14056), .I2(n14055), .O(n14058) );
  ND2DHD U15305 ( .I1(n9597), .I2(n14060), .O(n14061) );
  AN4CHD U15306 ( .I1(n14072), .I2(n14071), .I3(n6707), .I4(n14070), .O(n14073) );
  ND2DHD U15307 ( .I1(n8795), .I2(n14079), .O(n14089) );
  ND2DHD U15308 ( .I1(n14081), .I2(n6707), .O(n14086) );
  ND3CHD U15309 ( .I1(n6936), .I2(n14083), .I3(n14082), .O(n14085) );
  AOI22BHD U15310 ( .A1(n7017), .A2(KEY_88), .B1(n13292), .B2(n14094), .O(n14095) );
  OAI112BHD U15311 ( .C1(n10912), .C2(n14097), .A1(n14096), .B1(n14095), .O(n14099) );
  OAI22CHD U15312 ( .A1(n14880), .A2(n15513), .B1(n15512), .B2(n14608), .O(n14098) );
  AOI22BHD U15313 ( .A1(n15492), .A2(DIN_109), .B1(n7017), .B2(KEY_109), .O(n14105) );
  AOI22BHD U15314 ( .A1(n15492), .A2(DIN_45), .B1(n7017), .B2(KEY_45), .O(n14113) );
  AOI22BHD U15315 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _104), .B1(n15504), .B2(_i_CLEFIA128_keyK _40), .O(n14117) );
  AOI22BHD U15316 ( .A1(n7017), .A2(KEY_72), .B1(n13292), .B2(n14118), .O(n14119) );
  OAI112BHD U15317 ( .C1(n10912), .C2(n14121), .A1(n14120), .B1(n14119), .O(n14123) );
  OAI22CHD U15318 ( .A1(n15385), .A2(n15450), .B1(n15512), .B2(n15386), .O(n14122) );
  AOI22BHD U15319 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _96), .B1(n15504), .B2(_i_CLEFIA128_keyK _32), .O(n14127) );
  AOI22BHD U15320 ( .A1(n7017), .A2(KEY_64), .B1(n13292), .B2(n14128), .O(n14129) );
  OAI112BHD U15321 ( .C1(n10912), .C2(n14131), .A1(n14130), .B1(n14129), .O(n14133) );
  OAI22CHD U15322 ( .A1(n15511), .A2(n15513), .B1(n15512), .B2(n15514), .O(n14132) );
  NR2CHD U15323 ( .I1(n14133), .I2(n14132), .O(n14134) );
  AOI22BHD U15324 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _91), .B1(n15504), .B2(_i_CLEFIA128_keyK _27), .O(n14146) );
  AOI22BHD U15325 ( .A1(n7045), .A2(n14136), .B1(n15504), .B2(n14135), .O(n14145) );
  XNR2EHD U15326 ( .I1(n9013), .I2(n6847), .O(n14142) );
  AOI22BHD U15327 ( .A1(n7017), .A2(KEY_27), .B1(n13292), .B2(n14147), .O(n14148) );
  OAI112BHD U15328 ( .C1(n10912), .C2(n14150), .A1(n14149), .B1(n14148), .O(n14152) );
  OAI22CHD U15329 ( .A1(n14291), .A2(n15513), .B1(n15512), .B2(n15075), .O(n14151) );
  AOI22BHD U15330 ( .A1(n7045), .A2(n14155), .B1(n15504), .B2(n14154), .O(n14157) );
  XNR3EHD U15331 ( .I1(DOUT_81), .I2(n9775), .I3(n14351), .O(n14156) );
  XNR2KHD U15332 ( .I1(n14156), .I2(n14695), .O(n14575) );
  AOI22BHD U15333 ( .A1(n7017), .A2(KEY_81), .B1(n13292), .B2(n14158), .O(n14159) );
  OAI112BHD U15334 ( .C1(n10912), .C2(n14161), .A1(n14160), .B1(n14159), .O(n14163) );
  OAI22CHD U15335 ( .A1(n15141), .A2(n15513), .B1(n15512), .B2(n14871), .O(n14162) );
  AOI22BHD U15336 ( .A1(n15492), .A2(DIN_100), .B1(n7017), .B2(KEY_100), .O(n14165) );
  ND2DHD U15337 ( .I1(n9817), .I2(n15500), .O(n14174) );
  AOI22BHD U15338 ( .A1(n15492), .A2(DIN_117), .B1(n7017), .B2(KEY_117), .O(n14172) );
  AOI22BHD U15339 ( .A1(n15492), .A2(DIN_53), .B1(n7017), .B2(KEY_53), .O(n14176) );
  AOI22BHD U15340 ( .A1(n15492), .A2(DIN_36), .B1(n7017), .B2(KEY_36), .O(n14180) );
  OA12EHD U15341 ( .B1(n15499), .B2(n14983), .A1(n14180), .O(n14181) );
  AOI22BHD U15342 ( .A1(n7045), .A2(n14183), .B1(n15504), .B2(n14182), .O(n14185) );
  AOI22BHD U15343 ( .A1(n7017), .A2(KEY_93), .B1(n13292), .B2(n14186), .O(n14187) );
  OAI112BHD U15344 ( .C1(n10912), .C2(n14189), .A1(n14188), .B1(n14187), .O(n14191) );
  OAI22CHD U15345 ( .A1(n15159), .A2(n15450), .B1(n15512), .B2(n15160), .O(n14190) );
  ND2HHD U15346 ( .I1(n9779), .I2(n15500), .O(n14198) );
  AOI22BHD U15347 ( .A1(n15492), .A2(DIN_59), .B1(n7017), .B2(KEY_59), .O(n14195) );
  OA12EHD U15348 ( .B1(n15499), .B2(n15075), .A1(n14195), .O(n14196) );
  AOI22BHD U15349 ( .A1(n15492), .A2(DIN_123), .B1(n7017), .B2(KEY_123), .O(n14199) );
  OA12EHD U15350 ( .B1(n15499), .B2(n14291), .A1(n14199), .O(n14200) );
  AOI22BHD U15351 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _109), .B1(n15504), .B2(_i_CLEFIA128_keyK _45), .O(n14203) );
  AOI22BHD U15352 ( .A1(n7017), .A2(KEY_77), .B1(n13292), .B2(n14204), .O(n14205) );
  OAI112BHD U15353 ( .C1(n10912), .C2(n14207), .A1(n14206), .B1(n14205), .O(n14209) );
  OAI22CHD U15354 ( .A1(n15223), .A2(n15450), .B1(n15512), .B2(n15224), .O(n14208) );
  NR2CHD U15355 ( .I1(n14209), .I2(n14208), .O(n14210) );
  AOI22BHD U15356 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _101), .B1(n15504), .B2(_i_CLEFIA128_keyK _37), .O(n14217) );
  AOI22BHD U15357 ( .A1(n7045), .A2(n14212), .B1(n15504), .B2(n14211), .O(n14216) );
  AOI22BHD U15358 ( .A1(n7017), .A2(KEY_69), .B1(n13292), .B2(n14218), .O(n14219) );
  OAI112BHD U15359 ( .C1(n10912), .C2(n14221), .A1(n14220), .B1(n14219), .O(n14223) );
  OAI22CHD U15360 ( .A1(n15043), .A2(n15513), .B1(n15512), .B2(n15030), .O(n14222) );
  NR2CHD U15361 ( .I1(n14223), .I2(n14222), .O(n14224) );
  AOI22BHD U15362 ( .A1(n7045), .A2(n14226), .B1(n15504), .B2(n14225), .O(n14232) );
  AOI22BHD U15363 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _97), .B1(n15504), .B2(_i_CLEFIA128_keyK _33), .O(n14231) );
  XOR2EHD U15364 ( .I1(n14351), .I2(n14227), .O(n14230) );
  AOI22BHD U15365 ( .A1(n7017), .A2(KEY_65), .B1(n13292), .B2(n14233), .O(n14234) );
  OAI112BHD U15366 ( .C1(n10912), .C2(n14236), .A1(n14235), .B1(n14234), .O(n14238) );
  OAI22CHD U15367 ( .A1(n15258), .A2(n15513), .B1(n15512), .B2(n15271), .O(n14237) );
  AOI22BHD U15368 ( .A1(n7045), .A2(n14242), .B1(n15504), .B2(n14241), .O(n14248) );
  AOI22BHD U15369 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _69), .B1(n15504), .B2(_i_CLEFIA128_keyK _5), .O(n14247) );
  AOI22BHD U15370 ( .A1(n7017), .A2(KEY_5), .B1(n13292), .B2(n14249), .O(n14250) );
  OAI112BHD U15371 ( .C1(n10912), .C2(n14252), .A1(n14251), .B1(n14250), .O(n14254) );
  OAI22CHD U15372 ( .A1(n15030), .A2(n15450), .B1(n15512), .B2(n15043), .O(n14253) );
  AOI22BHD U15373 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _85), .B1(n15504), .B2(_i_CLEFIA128_keyK _21), .O(n14258) );
  AOI22BHD U15374 ( .A1(n7017), .A2(KEY_21), .B1(n13292), .B2(n14259), .O(n14260) );
  OAI112BHD U15375 ( .C1(n10912), .C2(n14262), .A1(n14261), .B1(n14260), .O(n14264) );
  OAI22CHD U15376 ( .A1(n14302), .A2(n15513), .B1(n15512), .B2(n14828), .O(n14263) );
  AOI22BHD U15377 ( .A1(n15492), .A2(DIN_44), .B1(n7017), .B2(KEY_44), .O(n14266) );
  OA12EHD U15378 ( .B1(n14633), .B2(n11129), .A1(n14267), .O(n14268) );
  AOI22BHD U15379 ( .A1(n15492), .A2(DIN_108), .B1(n7017), .B2(KEY_108), .O(n14270) );
  OA12EHD U15380 ( .B1(n14633), .B2(n15513), .A1(n14271), .O(n14272) );
  AOI22BHD U15381 ( .A1(n7017), .A2(KEY_92), .B1(n13292), .B2(n14277), .O(n14278) );
  OAI112BHD U15382 ( .C1(n10912), .C2(n14280), .A1(n14279), .B1(n14278), .O(n14282) );
  OAI22CHD U15383 ( .A1(n14924), .A2(n15513), .B1(n15512), .B2(n14321), .O(n14281) );
  AOI22BHD U15384 ( .A1(n7017), .A2(KEY_91), .B1(n13292), .B2(n14287), .O(n14288) );
  OAI112BHD U15385 ( .C1(n10912), .C2(n14290), .A1(n14289), .B1(n14288), .O(n14293) );
  OAI22CHD U15386 ( .A1(n15075), .A2(n15450), .B1(n15512), .B2(n14291), .O(n14292) );
  AOI22BHD U15387 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _117), .B1(n15504), .B2(_i_CLEFIA128_keyK _53), .O(n14297) );
  AOI22BHD U15388 ( .A1(n7017), .A2(KEY_85), .B1(n13292), .B2(n14298), .O(n14299) );
  OAI112BHD U15389 ( .C1(n10912), .C2(n14301), .A1(n14300), .B1(n14299), .O(n14304) );
  OAI22CHD U15390 ( .A1(n14828), .A2(n15513), .B1(n15512), .B2(n14302), .O(n14303) );
  AOI22BHD U15391 ( .A1(n7017), .A2(KEY_76), .B1(n13292), .B2(n14308), .O(n14309) );
  OAI112BHD U15392 ( .C1(n10912), .C2(n14311), .A1(n14310), .B1(n14309), .O(n14313) );
  OAI22CHD U15393 ( .A1(n15015), .A2(n15513), .B1(n15512), .B2(n15345), .O(n14312) );
  NR2CHD U15394 ( .I1(n14313), .I2(n14312), .O(n14314) );
  AOI22BHD U15395 ( .A1(n7017), .A2(KEY_28), .B1(n13292), .B2(n14317), .O(n14318) );
  OAI112BHD U15396 ( .C1(n10912), .C2(n14320), .A1(n14319), .B1(n14318), .O(n14323) );
  OAI22CHD U15397 ( .A1(n14321), .A2(n15450), .B1(n15512), .B2(n14924), .O(n14322) );
  XOR2EHD U15398 ( .I1(DOUT_67), .I2(n14327), .O(n14330) );
  AOI22BHD U15399 ( .A1(n7017), .A2(KEY_67), .B1(n13292), .B2(n14334), .O(n14335) );
  OAI112BHD U15400 ( .C1(n10912), .C2(n14337), .A1(n14336), .B1(n14335), .O(n14339) );
  OAI22CHD U15401 ( .A1(n15055), .A2(n15450), .B1(n15400), .B2(n15512), .O(n14338) );
  AOI22BHD U15402 ( .A1(n15492), .A2(DIN_116), .B1(n7017), .B2(KEY_116), .O(n14341) );
  AOI22BHD U15403 ( .A1(n15492), .A2(DIN_52), .B1(n7017), .B2(KEY_52), .O(n14346) );
  OAI12CHD U15404 ( .B1(n15499), .B2(n14384), .A1(n14346), .O(n14348) );
  AOI22BHD U15405 ( .A1(n7017), .A2(KEY_74), .B1(n13292), .B2(n14354), .O(n14355) );
  OAI112BHD U15406 ( .C1(n10912), .C2(n14357), .A1(n14356), .B1(n14355), .O(n14359) );
  OAI22CHD U15407 ( .A1(n14802), .A2(n15513), .B1(n15512), .B2(n15393), .O(n14358) );
  XNR3EHD U15408 ( .I1(n14365), .I2(n14364), .I3(n14363), .O(n14366) );
  AOI22BHD U15409 ( .A1(n7017), .A2(KEY_83), .B1(n13292), .B2(n14369), .O(n14370) );
  OAI112BHD U15410 ( .C1(n10912), .C2(n14372), .A1(n14371), .B1(n14370), .O(n14374) );
  OAI22CHD U15411 ( .A1(n15491), .A2(n15450), .B1(n15512), .B2(n15488), .O(n14373) );
  AOI22BHD U15412 ( .A1(n7017), .A2(KEY_84), .B1(n13292), .B2(n14379), .O(n14380) );
  OAI112BHD U15413 ( .C1(n10912), .C2(n14382), .A1(n14381), .B1(n14380), .O(n14386) );
  OAI22CHD U15414 ( .A1(n14384), .A2(n15513), .B1(n15512), .B2(n14383), .O(n14385) );
  AOI22BHD U15415 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _107), .B1(n15504), .B2(_i_CLEFIA128_keyK _43), .O(n14390) );
  AOI22BHD U15416 ( .A1(n7045), .A2(n11857), .B1(n15504), .B2(n14388), .O(n14389) );
  AOI22BHD U15417 ( .A1(n7017), .A2(KEY_75), .B1(n13292), .B2(n14391), .O(n14392) );
  OAI112BHD U15418 ( .C1(n10912), .C2(n14394), .A1(n14393), .B1(n14392), .O(n14396) );
  OAI22CHD U15419 ( .A1(n15316), .A2(n15513), .B1(n15512), .B2(n15317), .O(n14395) );
  NR2IHD U15420 ( .I1(_i_CLEFIA128_state_reg _1), .I2(_i_CLEFIA128_state_reg _0), .O(n14434) );
  ND2DHD U15421 ( .I1(n14401), .I2(n14683), .O(n14402) );
  ND2DHD U15422 ( .I1(n14402), .I2(n14430), .O(n14708) );
  OA22EHD U15423 ( .A1(n14685), .A2(n14688), .B1(n14721), .B2(n14719), .O(n14429) );
  NR2CHD U15424 ( .I1(n14429), .I2(n14404), .O(n14713) );
  AN2B1CHD U15425 ( .I1(n14709), .B1(n14713), .O(n14406) );
  ND2HHD U15426 ( .I1(n14407), .I2(n14434), .O(n14741) );
  ND2DHD U15427 ( .I1(n14410), .I2(n14409), .O(n14716) );
  NR2CHD U15428 ( .I1(n14414), .I2(n14420), .O(n14418) );
  MXL2CHD U15429 ( .A(n14417), .B(n14416), .S(n14415), .OB(n6372) );
  OAI22CHD U15430 ( .A1(_i_CLEFIA128_rndcnt_reg _3), .A2(n14420), .B1(n14709), .B2(n14419), .O(n14421) );
  NR2CHD U15431 ( .I1(n14716), .I2(n14421), .O(n14422) );
  AN2HHD U15432 ( .I1(n14425), .I2(n14434), .O(n14426) );
  NR2CHD U15433 ( .I1(SRST), .I2(n14426), .O(n15522) );
  NR2CHD U15434 ( .I1(n14427), .I2(n14426), .O(n14428) );
  ND2DHD U15435 ( .I1(n14429), .I2(n14428), .O(n14431) );
  MAOI1CHD U15436 ( .A1(n14433), .A2(_i_CLEFIA128_CON_T_x _2), .B1(n14432), .B2(n14753), .O(n14436) );
  AN2HHD U15437 ( .I1(n14432), .I2(n14434), .O(n14748) );
  ND3CHD U15438 ( .I1(n14437), .I2(n14436), .I3(n14468), .O(n6363) );
  MAOI1CHD U15439 ( .A1(n14433), .A2(_i_CLEFIA128_CON_T_x _8), .B1(n14432), .B2(n14736), .O(n14438) );
  ND2DHD U15440 ( .I1(n14748), .I2(n15492), .O(n14718) );
  ND3CHD U15441 ( .I1(n14439), .I2(n14438), .I3(n14718), .O(n6357) );
  ND2DHD U15442 ( .I1(n14433), .I2(_i_CLEFIA128_CON_T_x _0), .O(n14743) );
  ND3CHD U15443 ( .I1(n14442), .I2(n14441), .I3(n14741), .O(n6365) );
  ND2DHD U15444 ( .I1(n14433), .I2(n14443), .O(n14742) );
  ND3CHD U15445 ( .I1(n14453), .I2(n14452), .I3(n14451), .O(n6352) );
  ND3CHD U15446 ( .I1(n14458), .I2(n14457), .I3(n14456), .O(n6360) );
  ND3CHD U15447 ( .I1(n14463), .I2(n14462), .I3(n14461), .O(n6354) );
  AOI22BHD U15448 ( .A1(_i_CLEFIA128_CON_T_xi _11), .A2(n14475), .B1(n14433), .B2(_i_CLEFIA128_CON_T_x _12), .O(n14466) );
  ND2DHD U15449 ( .I1(n14467), .I2(n14466), .O(n6353) );
  MAOI1CHD U15450 ( .A1(n14433), .A2(_i_CLEFIA128_CON_T_x _14), .B1(n14432), .B2(n14469), .O(n14470) );
  ND3CHD U15451 ( .I1(n14471), .I2(n14473), .I3(n14470), .O(n6351) );
  AOI22BHD U15452 ( .A1(n14433), .A2(_i_CLEFIA128_CON_T_x _3), .B1(n14475), .B2(_i_CLEFIA128_CON_T_xi_2 ), .O(n14472) );
  ND3CHD U15453 ( .I1(n14474), .I2(n14473), .I3(n14472), .O(n6362) );
  AOI22BHD U15454 ( .A1(n14433), .A2(_i_CLEFIA128_CON_T_x _10), .B1(n14475), .B2(_i_CLEFIA128_CON_T_xi _9), .O(n14476) );
  ND3CHD U15455 ( .I1(n14477), .I2(n14476), .I3(n14741), .O(n6355) );
  OAI112BHD U15456 ( .C1(n15422), .C2(n15352), .A1(n14479), .B1(n14478), .O(n14480) );
  OAI112BHD U15457 ( .C1(n15422), .C2(n14556), .A1(n14485), .B1(n14484), .O(n14486) );
  OAI12CHD U15458 ( .B1(n14615), .B2(n15416), .A1(n14488), .O(n6324) );
  OAI112BHD U15459 ( .C1(n15422), .C2(n15398), .A1(n14495), .B1(n14494), .O(n14496) );
  OAI12CHD U15460 ( .B1(n15486), .B2(n15416), .A1(n14498), .O(n6341) );
  OAI112BHD U15461 ( .C1(n15422), .C2(n14988), .A1(n14501), .B1(n14500), .O(n14502) );
  OAI12CHD U15462 ( .B1(n14573), .B2(n15416), .A1(n14504), .O(n6331) );
  OAI112BHD U15463 ( .C1(n15422), .C2(n15035), .A1(n14506), .B1(n14505), .O(n14507) );
  OAI12CHD U15464 ( .B1(n15374), .B2(n15416), .A1(n14509), .O(n6332) );
  OAI112BHD U15465 ( .C1(n15422), .C2(n15096), .A1(n14511), .B1(n14510), .O(n14512) );
  OAI12CHD U15466 ( .B1(n9697), .B2(n15416), .A1(n14514), .O(n6279) );
  OAI112BHD U15467 ( .C1(n15422), .C2(n15046), .A1(n14516), .B1(n14515), .O(n14517) );
  OAI12CHD U15468 ( .B1(n15503), .B2(n15416), .A1(n14519), .O(n6319) );
  OAI112BHD U15469 ( .C1(n15422), .C2(n14975), .A1(n14521), .B1(n14520), .O(n14522) );
  OAI12CHD U15470 ( .B1(n14525), .B2(n15416), .A1(n14524), .O(n6318) );
  OAI112BHD U15471 ( .C1(n15422), .C2(n15407), .A1(n14527), .B1(n14526), .O(n14528) );
  NR2CHD U15472 ( .I1(n14529), .I2(n14528), .O(n14530) );
  OAI112BHD U15473 ( .C1(n15422), .C2(n8902), .A1(n14532), .B1(n14531), .O(n14533) );
  OAI12CHD U15474 ( .B1(n15377), .B2(n15416), .A1(n14535), .O(n6269) );
  OAI112BHD U15475 ( .C1(n15422), .C2(n15029), .A1(n14537), .B1(n14536), .O(n14538) );
  OAI12CHD U15476 ( .B1(n7082), .B2(n15416), .A1(n14540), .O(n6346) );
  OAI112BHD U15477 ( .C1(n15422), .C2(n15040), .A1(n14542), .B1(n14541), .O(n14543) );
  OAI112BHD U15478 ( .C1(n15422), .C2(n14972), .A1(n14547), .B1(n14546), .O(n14548) );
  OAI12CHD U15479 ( .B1(n14613), .B2(n15416), .A1(n14550), .O(n6261) );
  OAI112BHD U15480 ( .C1(n15422), .C2(n15409), .A1(n14552), .B1(n14551), .O(n14553) );
  OAI12CHD U15481 ( .B1(n15449), .B2(n15416), .A1(n14555), .O(n6271) );
  OAI112BHD U15482 ( .C1(n15422), .C2(n14979), .A1(n14559), .B1(n14558), .O(n14560) );
  OAI12CHD U15483 ( .B1(n9089), .B2(n15416), .A1(n14562), .O(n6254) );
  AOI22BHD U15484 ( .A1(n15492), .A2(DIN_113), .B1(n7017), .B2(KEY_113), .O(n14563) );
  OA12EHD U15485 ( .B1(n15499), .B2(n14871), .A1(n14563), .O(n14564) );
  OAI12CHD U15486 ( .B1(n14575), .B2(n15513), .A1(n14565), .O(n6207) );
  OAI112BHD U15487 ( .C1(n15422), .C2(n15069), .A1(n14567), .B1(n14566), .O(n14568) );
  OAI12CHD U15488 ( .B1(n14575), .B2(n15416), .A1(n14570), .O(n6268) );
  AOI22BHD U15489 ( .A1(n15492), .A2(DIN_49), .B1(n7017), .B2(KEY_49), .O(n14571) );
  OA12EHD U15490 ( .B1(n14573), .B2(n15450), .A1(n14572), .O(n14574) );
  OAI12CHD U15491 ( .B1(n14575), .B2(n11129), .A1(n14574), .O(n6175) );
  OAI112BHD U15492 ( .C1(n15422), .C2(n15172), .A1(n14577), .B1(n14576), .O(n14578) );
  OAI12CHD U15493 ( .B1(n10008), .B2(n15416), .A1(n14580), .O(n6256) );
  OAI112BHD U15494 ( .C1(n15422), .C2(n15194), .A1(n14582), .B1(n14581), .O(n14583) );
  OAI112BHD U15495 ( .C1(n15422), .C2(n15257), .A1(n14587), .B1(n14586), .O(n14588) );
  OAI12CHD U15496 ( .B1(n7613), .B2(n15416), .A1(n14590), .O(n6343) );
  OAI112BHD U15497 ( .C1(n15422), .C2(n15300), .A1(n14592), .B1(n14591), .O(n14593) );
  OAI112BHD U15498 ( .C1(n15422), .C2(n15399), .A1(n14597), .B1(n14596), .O(n14598) );
  OAI12CHD U15499 ( .B1(n14601), .B2(n15416), .A1(n14600), .O(n6257) );
  OAI112BHD U15500 ( .C1(n15422), .C2(n15244), .A1(n14603), .B1(n14602), .O(n14604) );
  AOI22BHD U15501 ( .A1(n15492), .A2(DIN_120), .B1(n7017), .B2(KEY_120), .O(n14607) );
  OA12EHD U15502 ( .B1(n14613), .B2(n15513), .A1(n14609), .O(n14610) );
  OAI12CHD U15503 ( .B1(n14615), .B2(n11129), .A1(n14610), .O(n6214) );
  AOI22BHD U15504 ( .A1(n15492), .A2(DIN_56), .B1(n7017), .B2(KEY_56), .O(n14611) );
  OA12EHD U15505 ( .B1(n15499), .B2(n14880), .A1(n14611), .O(n14612) );
  OA12EHD U15506 ( .B1(n14613), .B2(n15512), .A1(n14612), .O(n14614) );
  OAI12CHD U15507 ( .B1(n14615), .B2(n15513), .A1(n14614), .O(n6182) );
  OAI112BHD U15508 ( .C1(n15422), .C2(n15128), .A1(n14617), .B1(n14616), .O(n14618) );
  OAI12CHD U15509 ( .B1(n14621), .B2(n15416), .A1(n14620), .O(n6258) );
  OAI112BHD U15510 ( .C1(n15422), .C2(n14919), .A1(n14623), .B1(n14622), .O(n14624) );
  OAI12CHD U15511 ( .B1(n15134), .B2(n15416), .A1(n14626), .O(n6267) );
  AOI22BHD U15512 ( .A1(n15492), .A2(DIN_50), .B1(n7017), .B2(KEY_50), .O(n14627) );
  OAI112BHD U15513 ( .C1(n15422), .C2(n15061), .A1(n14629), .B1(n14628), .O(n14630) );
  OAI112BHD U15514 ( .C1(n15422), .C2(n15344), .A1(n14638), .B1(n14637), .O(n14639) );
  OAI12CHD U15515 ( .B1(n6904), .B2(n15416), .A1(n14641), .O(n6283) );
  AOI22BHD U15516 ( .A1(n15492), .A2(DIN_34), .B1(n7017), .B2(KEY_34), .O(n14642) );
  OA12EHD U15517 ( .B1(n14647), .B2(n15513), .A1(n14643), .O(n14644) );
  OAI12CHD U15518 ( .B1(n6904), .B2(n11129), .A1(n14644), .O(n6160) );
  AOI22BHD U15519 ( .A1(n15492), .A2(DIN_98), .B1(n7017), .B2(KEY_98), .O(n14645) );
  OA12EHD U15520 ( .B1(n15499), .B2(n15329), .A1(n14645), .O(n14646) );
  OAI12CHD U15521 ( .B1(n6904), .B2(n15513), .A1(n14648), .O(n6192) );
  OAI112BHD U15522 ( .C1(n15422), .C2(n15263), .A1(n14650), .B1(n14649), .O(n14651) );
  OAI12CHD U15523 ( .B1(n7970), .B2(n15416), .A1(n14653), .O(n6329) );
  OAI112BHD U15524 ( .C1(n15422), .C2(n15298), .A1(n14655), .B1(n14654), .O(n14656) );
  NR2CHD U15525 ( .I1(n14657), .I2(n14656), .O(n14658) );
  OAI112BHD U15526 ( .C1(n15422), .C2(n15293), .A1(n14660), .B1(n14659), .O(n14661) );
  OAI112BHD U15527 ( .C1(n15422), .C2(n15089), .A1(n14665), .B1(n14664), .O(n14666) );
  AOI22BHD U15528 ( .A1(n15492), .A2(DIN_37), .B1(n7017), .B2(KEY_37), .O(n14669) );
  AOI22BHD U15529 ( .A1(n15492), .A2(DIN_101), .B1(n7017), .B2(KEY_101), .O(n14670) );
  OA12EHD U15530 ( .B1(n15499), .B2(n15030), .A1(n14670), .O(n14671) );
  AOI22BHD U15531 ( .A1(n15492), .A2(DIN_99), .B1(n7017), .B2(KEY_99), .O(n14672) );
  AOI22BHD U15532 ( .A1(n15492), .A2(DIN_35), .B1(n7017), .B2(KEY_35), .O(n14675) );
  ND3CHD U15533 ( .I1(n14688), .I2(n14680), .I3(n14679), .O(n14681) );
  MXL2CHD U15534 ( .A(n14692), .B(n14691), .S(n14695), .OB(n14706) );
  ND2DHD U15535 ( .I1(n14695), .I2(n14692), .O(n14693) );
  OAI12CHD U15536 ( .B1(n14695), .B2(n14694), .A1(n14693), .O(n14696) );
  AOI22BHD U15537 ( .A1(n7017), .A2(KEY_90), .B1(n13292), .B2(n14697), .O(n14698) );
  OAI112BHD U15538 ( .C1(n10912), .C2(n14700), .A1(n14699), .B1(n14698), .O(n14702) );
  OAI22CHD U15539 ( .A1(n14959), .A2(n15513), .B1(n15512), .B2(n15337), .O(n14701) );
  OAI112BHD U15540 ( .C1(n9538), .C2(n14706), .A1(n14704), .B1(n14703), .O(n6132) );
  NR2CHD U15541 ( .I1(n8189), .I2(n7048), .O(n14710) );
  ND2DHD U15542 ( .I1(n14712), .I2(n14711), .O(n6370) );
  ND3CHD U15543 ( .I1(n14723), .I2(_i_CLEFIA128_state_reg _1), .I3(n15522), .O(n14717) );
  ND3CHD U15544 ( .I1(n14741), .I2(n14725), .I3(n14724), .O(n6368) );
  OAI112BHD U15545 ( .C1(n14731), .C2(n14752), .A1(n14730), .B1(n14729), .O(n6356) );
  OAI112BHD U15546 ( .C1(n14736), .C2(n14752), .A1(n14735), .B1(n14734), .O(n6358) );
  ND2DHD U15547 ( .I1(n14746), .I2(n14745), .O(n6361) );
  OAI112BHD U15548 ( .C1(n14753), .C2(n14752), .A1(n14751), .B1(n14750), .O(n6364) );
  AOI22BHD U15549 ( .A1(n7045), .A2(n14755), .B1(n15504), .B2(n14754), .O(n14765) );
  AO22CHD U15550 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _127), .B1(n15504), .B2(_i_CLEFIA128_keyK _63), .O(n14756) );
  ND2DHD U15551 ( .I1(n14766), .I2(n14756), .O(n14764) );
  AOI22BHD U15552 ( .A1(n7017), .A2(KEY_95), .B1(n13292), .B2(n14757), .O(n14758) );
  OAI112BHD U15553 ( .C1(n10912), .C2(n14760), .A1(n14759), .B1(n14758), .O(n14762) );
  OAI22CHD U15554 ( .A1(n14866), .A2(n15513), .B1(n15512), .B2(n15417), .O(n14761) );
  OAI112BHD U15555 ( .C1(n9089), .C2(n14765), .A1(n14764), .B1(n14763), .O(n6127) );
  AOI22BHD U15556 ( .A1(n15492), .A2(DIN_39), .B1(n7017), .B2(KEY_39), .O(n14769) );
  OAI112BHD U15557 ( .C1(n15486), .C2(n15513), .A1(n14771), .B1(n14770), .O(n6165) );
  AOI22BHD U15558 ( .A1(n7045), .A2(n14773), .B1(n15504), .B2(n14772), .O(n14783) );
  AO22CHD U15559 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _71), .B1(n15504), .B2(_i_CLEFIA128_keyK _7), .O(n14774) );
  AOI22BHD U15560 ( .A1(n7017), .A2(KEY_7), .B1(n13292), .B2(n14775), .O(n14776) );
  OAI112BHD U15561 ( .C1(n10912), .C2(n14778), .A1(n14777), .B1(n14776), .O(n14780) );
  OAI22CHD U15562 ( .A1(n15483), .A2(n15513), .B1(n15512), .B2(n15475), .O(n14779) );
  OAI112BHD U15563 ( .C1(n15486), .C2(n14783), .A1(n14782), .B1(n14781), .O(n6120) );
  AOI22BHD U15564 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _79), .B1(n15504), .B2(_i_CLEFIA128_keyK _15), .O(n14795) );
  AO22CHD U15565 ( .A1(n7045), .A2(n14785), .B1(n15504), .B2(n14784), .O(n14786) );
  AOI22BHD U15566 ( .A1(n7017), .A2(KEY_15), .B1(n13292), .B2(n14787), .O(n14788) );
  OAI112BHD U15567 ( .C1(n10912), .C2(n14790), .A1(n14789), .B1(n14788), .O(n14792) );
  OAI22CHD U15568 ( .A1(n15360), .A2(n15513), .B1(n15512), .B2(n15361), .O(n14791) );
  OAI112BHD U15569 ( .C1(n15207), .C2(n14795), .A1(n14794), .B1(n14793), .O(n6112) );
  OAI12CHD U15570 ( .B1(n13277), .B2(n15046), .A1(n14799), .O(n14800) );
  AOI22BHD U15571 ( .A1(n15492), .A2(DIN_42), .B1(n7017), .B2(KEY_42), .O(n14801) );
  AOI22BHD U15572 ( .A1(n15492), .A2(DIN_125), .B1(n7017), .B2(KEY_125), .O(n14806) );
  AOI22BHD U15573 ( .A1(n15492), .A2(DIN_61), .B1(n7017), .B2(KEY_61), .O(n14807) );
  OAI12CHD U15574 ( .B1(n13277), .B2(n14817), .A1(n14811), .O(n14812) );
  OAI112BHD U15575 ( .C1(n13277), .C2(n15208), .A1(n14819), .B1(n14818), .O(n6249) );
  OAI112BHD U15576 ( .C1(n13277), .C2(n15236), .A1(n14823), .B1(n14822), .O(n6315) );
  OAI112BHD U15577 ( .C1(n13277), .C2(n14945), .A1(n14827), .B1(n14826), .O(n6310) );
  OAI112BHD U15578 ( .C1(n13277), .C2(n14919), .A1(n14832), .B1(n14831), .O(n6296) );
  OAI112BHD U15579 ( .C1(n13277), .C2(n14939), .A1(n14845), .B1(n14844), .O(n6239) );
  OAI12CHD U15580 ( .B1(n13277), .B2(n7392), .A1(n14848), .O(n14849) );
  OAI112BHD U15581 ( .C1(n13277), .C2(n14953), .A1(n14853), .B1(n14852), .O(n6253) );
  OAI112BHD U15582 ( .C1(n13277), .C2(n15061), .A1(n14857), .B1(n14856), .O(n6288) );
  OAI112BHD U15583 ( .C1(n13277), .C2(n14864), .A1(n14861), .B1(n14860), .O(n6238) );
  OAI112BHD U15584 ( .C1(n13277), .C2(n15409), .A1(n14870), .B1(n14869), .O(n6286) );
  OAI112BHD U15585 ( .C1(n13277), .C2(n15146), .A1(n14875), .B1(n14874), .O(n6236) );
  OAI12CHD U15586 ( .B1(n13277), .B2(n15140), .A1(n14878), .O(n14879) );
  OAI112BHD U15587 ( .C1(n13277), .C2(n15296), .A1(n14884), .B1(n14883), .O(n6293) );
  AOI22BHD U15588 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _121), .B1(n15504), .B2(_i_CLEFIA128_keyK _57), .O(n14895) );
  AO22CHD U15589 ( .A1(n7045), .A2(n8081), .B1(n15504), .B2(n14885), .O(n14886) );
  AOI22BHD U15590 ( .A1(n7017), .A2(KEY_89), .B1(n13292), .B2(n14887), .O(n14888) );
  OAI112BHD U15591 ( .C1(n10912), .C2(n14890), .A1(n14889), .B1(n14888), .O(n14892) );
  OAI22CHD U15592 ( .A1(n15461), .A2(n15513), .B1(n15512), .B2(n15462), .O(n14891) );
  OAI112BHD U15593 ( .C1(n14913), .C2(n14895), .A1(n14894), .B1(n14893), .O(n6133) );
  OAI12CHD U15594 ( .B1(n13277), .B2(n15182), .A1(n14898), .O(n14899) );
  OAI112BHD U15595 ( .C1(n13277), .C2(n15194), .A1(n14903), .B1(n14902), .O(n6228) );
  OAI112BHD U15596 ( .C1(n13277), .C2(n15186), .A1(n14908), .B1(n14907), .O(n6299) );
  OAI12CHD U15597 ( .B1(n13277), .B2(n14954), .A1(n14911), .O(n14912) );
  OAI112BHD U15598 ( .C1(n13277), .C2(n14918), .A1(n14917), .B1(n14916), .O(n6303) );
  OAI112BHD U15599 ( .C1(n13277), .C2(n14930), .A1(n14929), .B1(n14928), .O(n6289) );
  OAI12CHD U15600 ( .B1(n13277), .B2(n14936), .A1(n14935), .O(n14937) );
  OAI12CHD U15601 ( .B1(n13277), .B2(n14943), .A1(n14942), .O(n14944) );
  OAI112BHD U15602 ( .C1(n13277), .C2(n14950), .A1(n14949), .B1(n14948), .O(n6246) );
  OAI112BHD U15603 ( .C1(n13277), .C2(n14957), .A1(n14956), .B1(n14955), .O(n6317) );
  AOI22BHD U15604 ( .A1(n15492), .A2(DIN_58), .B1(n7017), .B2(KEY_58), .O(n14958) );
  OAI12CHD U15605 ( .B1(n15499), .B2(n14959), .A1(n14958), .O(n14960) );
  OAI112BHD U15606 ( .C1(n13277), .C2(n15270), .A1(n14967), .B1(n14966), .O(n6302) );
  OAI112BHD U15607 ( .C1(n13277), .C2(n14972), .A1(n14971), .B1(n14970), .O(n6304) );
  OAI112BHD U15608 ( .C1(n13277), .C2(n14979), .A1(n14978), .B1(n14977), .O(n6311) );
  AOI22BHD U15609 ( .A1(n15492), .A2(DIN_97), .B1(n7017), .B2(KEY_97), .O(n14980) );
  OAI112BHD U15610 ( .C1(n15054), .C2(n15513), .A1(n14982), .B1(n14981), .O(n6191) );
  OAI112BHD U15611 ( .C1(n13277), .C2(n15172), .A1(n14987), .B1(n14986), .O(n6313) );
  XOR2EHD U15612 ( .I1(DOUT_73), .I2(n9923), .O(n14995) );
  ND2DHD U15613 ( .I1(n15024), .I2(n15500), .O(n14999) );
  AOI22BHD U15614 ( .A1(n15492), .A2(DIN_105), .B1(n7017), .B2(KEY_105), .O(n14997) );
  AOI22BHD U15615 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _105), .B1(n15504), .B2(_i_CLEFIA128_keyK _41), .O(n15011) );
  AO22CHD U15616 ( .A1(n7045), .A2(n15001), .B1(n15504), .B2(n15000), .O(n15002) );
  AOI22BHD U15617 ( .A1(n7017), .A2(KEY_73), .B1(n13292), .B2(n15003), .O(n15004) );
  OAI112BHD U15618 ( .C1(n10912), .C2(n15006), .A1(n15005), .B1(n15004), .O(n15008) );
  OAI22CHD U15619 ( .A1(n15115), .A2(n15513), .B1(n15512), .B2(n15106), .O(n15007) );
  OAI112BHD U15620 ( .C1(n15024), .C2(n15011), .A1(n15010), .B1(n15009), .O(n6149) );
  AOI22BHD U15621 ( .A1(n15492), .A2(DIN_41), .B1(n7017), .B2(KEY_41), .O(n15012) );
  OAI112BHD U15622 ( .C1(n13277), .C2(n15036), .A1(n15019), .B1(n15018), .O(n6305) );
  OAI12CHD U15623 ( .B1(n13277), .B2(n15042), .A1(n15022), .O(n15023) );
  OAI112BHD U15624 ( .C1(n13277), .C2(n15029), .A1(n15028), .B1(n15027), .O(n6234) );
  OAI112BHD U15625 ( .C1(n13277), .C2(n15035), .A1(n15034), .B1(n15033), .O(n6248) );
  OAI12CHD U15626 ( .B1(n13277), .B2(n15040), .A1(n15039), .O(n15041) );
  OAI112BHD U15627 ( .C1(n13277), .C2(n15050), .A1(n15049), .B1(n15048), .O(n6312) );
  ND2DHD U15628 ( .I1(n15200), .I2(n15500), .O(n15053) );
  AOI22BHD U15629 ( .A1(n15492), .A2(DIN_33), .B1(n7017), .B2(KEY_33), .O(n15051) );
  OAI112BHD U15630 ( .C1(n15054), .C2(n11129), .A1(n15053), .B1(n15052), .O(n6159) );
  OAI112BHD U15631 ( .C1(n13277), .C2(n15403), .A1(n15060), .B1(n15059), .O(n6314) );
  OAI12CHD U15632 ( .B1(n13277), .B2(n15290), .A1(n15065), .O(n15066) );
  AOI22BHD U15633 ( .A1(n15492), .A2(DIN_106), .B1(n7017), .B2(KEY_106), .O(n15068) );
  OAI112BHD U15634 ( .C1(n13277), .C2(n15301), .A1(n15080), .B1(n15079), .O(n6290) );
  OAI112BHD U15635 ( .C1(n13277), .C2(n15096), .A1(n15084), .B1(n15083), .O(n6223) );
  OAI112BHD U15636 ( .C1(n13277), .C2(n15092), .A1(n15088), .B1(n15087), .O(n6287) );
  OAI12CHD U15637 ( .B1(n13277), .B2(n15100), .A1(n15099), .O(n15101) );
  OAI112BHD U15638 ( .C1(n13277), .C2(n9474), .A1(n15105), .B1(n15104), .O(n6230) );
  OAI112BHD U15639 ( .C1(n13277), .C2(n15244), .A1(n15110), .B1(n15109), .O(n6244) );
  OAI112BHD U15640 ( .C1(n13277), .C2(n15247), .A1(n15114), .B1(n15113), .O(n6251) );
  OAI112BHD U15641 ( .C1(n13277), .C2(n15120), .A1(n15119), .B1(n15118), .O(n6308) );
  OAI112BHD U15642 ( .C1(n13277), .C2(n15128), .A1(n15127), .B1(n15126), .O(n6301) );
  AOI22BHD U15643 ( .A1(n15492), .A2(DIN_114), .B1(n7017), .B2(KEY_114), .O(n15129) );
  ND2DHD U15644 ( .I1(n15131), .I2(n11130), .O(n15132) );
  OAI112BHD U15645 ( .C1(n15134), .C2(n15513), .A1(n15133), .B1(n15132), .O(n6208) );
  OAI112BHD U15646 ( .C1(n13277), .C2(n15399), .A1(n15145), .B1(n15144), .O(n6300) );
  OAI12CHD U15647 ( .B1(n13277), .B2(n15150), .A1(n15149), .O(n15151) );
  AOI22BHD U15648 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _93), .B1(n15504), .B2(_i_CLEFIA128_keyK _29), .O(n15165) );
  AO22CHD U15649 ( .A1(n7045), .A2(n8173), .B1(n15504), .B2(n15153), .O(n15154) );
  AOI22BHD U15650 ( .A1(n7017), .A2(KEY_29), .B1(n13292), .B2(n15155), .O(n15156) );
  OAI112BHD U15651 ( .C1(n10912), .C2(n15158), .A1(n15157), .B1(n15156), .O(n15162) );
  OAI22CHD U15652 ( .A1(n15160), .A2(n15513), .B1(n15512), .B2(n15159), .O(n15161) );
  NR2CHD U15653 ( .I1(n15162), .I2(n15161), .O(n15163) );
  OAI112BHD U15654 ( .C1(n15171), .C2(n15165), .A1(n15164), .B1(n15163), .O(n6098) );
  OAI12CHD U15655 ( .B1(n13277), .B2(n15169), .A1(n15168), .O(n15170) );
  OAI12CHD U15656 ( .B1(n13277), .B2(n15176), .A1(n15175), .O(n15177) );
  OAI112BHD U15657 ( .C1(n13277), .C2(n15185), .A1(n15184), .B1(n15183), .O(n6306) );
  OAI12CHD U15658 ( .B1(n13277), .B2(n15191), .A1(n15190), .O(n15192) );
  OAI12CHD U15659 ( .B1(n13277), .B2(n15198), .A1(n15197), .O(n15199) );
  OAI12CHD U15660 ( .B1(n13277), .B2(n15205), .A1(n15204), .O(n15206) );
  OAI12CHD U15661 ( .B1(n13277), .B2(n15214), .A1(n15213), .O(n15215) );
  AOI22BHD U15662 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _77), .B1(n15504), .B2(_i_CLEFIA128_keyK _13), .O(n15229) );
  AOI22BHD U15663 ( .A1(n7017), .A2(KEY_13), .B1(n13292), .B2(n15219), .O(n15220) );
  OAI112BHD U15664 ( .C1(n10912), .C2(n15222), .A1(n15221), .B1(n15220), .O(n15226) );
  OAI22CHD U15665 ( .A1(n15224), .A2(n15513), .B1(n15512), .B2(n15223), .O(n15225) );
  OAI112BHD U15666 ( .C1(n15235), .C2(n15229), .A1(n15228), .B1(n15227), .O(n6114) );
  OAI12CHD U15667 ( .B1(n13277), .B2(n15233), .A1(n15232), .O(n15234) );
  OAI112BHD U15668 ( .C1(n13277), .C2(n15242), .A1(n15241), .B1(n15240), .O(n6237) );
  OAI112BHD U15669 ( .C1(n13277), .C2(n15257), .A1(n15256), .B1(n15255), .O(n6231) );
  OAI112BHD U15670 ( .C1(n13277), .C2(n15274), .A1(n15262), .B1(n15261), .O(n6316) );
  OAI12CHD U15671 ( .B1(n13277), .B2(n15267), .A1(n15266), .O(n15268) );
  OAI112BHD U15672 ( .C1(n13277), .C2(n15277), .A1(n15276), .B1(n15275), .O(n6252) );
  OAI112BHD U15673 ( .C1(n13277), .C2(n15284), .A1(n15283), .B1(n15282), .O(n6309) );
  OAI112BHD U15674 ( .C1(n13277), .C2(n15293), .A1(n15292), .B1(n15291), .O(n6295) );
  OAI12CHD U15675 ( .B1(n13277), .B2(n15298), .A1(n15297), .O(n15299) );
  AOI22BHD U15676 ( .A1(n15492), .A2(DIN_43), .B1(n7017), .B2(KEY_43), .O(n15308) );
  AOI22BHD U15677 ( .A1(n7017), .A2(KEY_11), .B1(n13292), .B2(n15312), .O(n15313) );
  OAI112BHD U15678 ( .C1(n10912), .C2(n15315), .A1(n15314), .B1(n15313), .O(n15319) );
  OAI22CHD U15679 ( .A1(n15317), .A2(n15513), .B1(n15512), .B2(n15316), .O(n15318) );
  AO22CHD U15680 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _98), .B1(n15504), .B2(_i_CLEFIA128_keyK _34), .O(n15324) );
  AOI22BHD U15681 ( .A1(n7017), .A2(KEY_66), .B1(n13292), .B2(n15325), .O(n15326) );
  OAI112BHD U15682 ( .C1(n10912), .C2(n15328), .A1(n15327), .B1(n15326), .O(n15332) );
  OAI22CHD U15683 ( .A1(n15330), .A2(n15513), .B1(n15512), .B2(n15329), .O(n15331) );
  OAI112BHD U15684 ( .C1(n13277), .C2(n15344), .A1(n15343), .B1(n15342), .O(n6227) );
  OAI112BHD U15685 ( .C1(n13277), .C2(n15352), .A1(n15351), .B1(n15350), .O(n6241) );
  AOI22BHD U15686 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _111), .B1(n15504), .B2(_i_CLEFIA128_keyK _47), .O(n15366) );
  AO22CHD U15687 ( .A1(n7045), .A2(n15354), .B1(n15504), .B2(n15353), .O(n15355) );
  AOI22BHD U15688 ( .A1(n7017), .A2(KEY_79), .B1(n13292), .B2(n15356), .O(n15357) );
  OAI112BHD U15689 ( .C1(n10912), .C2(n15359), .A1(n15358), .B1(n15357), .O(n15363) );
  OAI22CHD U15690 ( .A1(n15361), .A2(n15513), .B1(n15512), .B2(n15360), .O(n15362) );
  OAI112BHD U15691 ( .C1(n15367), .C2(n15366), .A1(n15365), .B1(n15364), .O(n6143) );
  AOI22BHD U15692 ( .A1(n15492), .A2(DIN_112), .B1(n7017), .B2(KEY_112), .O(n15368) );
  AOI22BHD U15693 ( .A1(n15492), .A2(DIN_48), .B1(n7017), .B2(KEY_48), .O(n15372) );
  OR2EHD U15694 ( .I1(n15513), .I2(n15374), .O(n15375) );
  OAI112BHD U15695 ( .C1(n15377), .C2(n11129), .A1(n15376), .B1(n15375), .O(n6174) );
  AOI22BHD U15696 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _72), .B1(n15504), .B2(_i_CLEFIA128_keyK _8), .O(n15391) );
  AO22CHD U15697 ( .A1(n7045), .A2(n15379), .B1(n15504), .B2(n15378), .O(n15380) );
  AOI22BHD U15698 ( .A1(n7017), .A2(KEY_8), .B1(n13292), .B2(n15381), .O(n15382) );
  OAI112BHD U15699 ( .C1(n10912), .C2(n15384), .A1(n15383), .B1(n15382), .O(n15388) );
  OAI22CHD U15700 ( .A1(n15386), .A2(n15513), .B1(n15512), .B2(n15385), .O(n15387) );
  OAI112BHD U15701 ( .C1(n15392), .C2(n15391), .A1(n15390), .B1(n15389), .O(n6119) );
  OAI112BHD U15702 ( .C1(n13277), .C2(n15398), .A1(n15397), .B1(n15396), .O(n6243) );
  OAI112BHD U15703 ( .C1(n13277), .C2(n15407), .A1(n15406), .B1(n15405), .O(n6250) );
  OAI12CHD U15704 ( .B1(n13277), .B2(n15413), .A1(n15412), .O(n15414) );
  OAI112BHD U15705 ( .C1(n13277), .C2(n15426), .A1(n15425), .B1(n15424), .O(n6222) );
  AOI22BHD U15706 ( .A1(n15492), .A2(DIN_102), .B1(n7017), .B2(KEY_102), .O(n15427) );
  OAI112BHD U15707 ( .C1(n9697), .C2(n15513), .A1(n15430), .B1(n15429), .O(n6196) );
  AOI22BHD U15708 ( .A1(n15492), .A2(DIN_55), .B1(n7017), .B2(KEY_55), .O(n15431) );
  OAI112BHD U15709 ( .C1(n6604), .C2(n15513), .A1(n15434), .B1(n15433), .O(n6181) );
  AOI22BHD U15710 ( .A1(n15492), .A2(DIN_119), .B1(n7017), .B2(KEY_119), .O(n15436) );
  AOI22BHD U15711 ( .A1(n15492), .A2(DIN_38), .B1(n7017), .B2(KEY_38), .O(n15441) );
  OAI112BHD U15712 ( .C1(n9697), .C2(n11129), .A1(n15444), .B1(n15443), .O(n6164) );
  AOI22BHD U15713 ( .A1(n15492), .A2(DIN_46), .B1(n7017), .B2(KEY_46), .O(n15445) );
  OA12EHD U15714 ( .B1(n15499), .B2(n15446), .A1(n15445), .O(n15447) );
  AOI22BHD U15715 ( .A1(n15492), .A2(DIN_110), .B1(n7017), .B2(KEY_110), .O(n15451) );
  OA12EHD U15716 ( .B1(n15499), .B2(n15452), .A1(n15451), .O(n15453) );
  AOI22BHD U15717 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _89), .B1(n15504), .B2(_i_CLEFIA128_keyK _25), .O(n15467) );
  AO22CHD U15718 ( .A1(n7045), .A2(n8051), .B1(n15504), .B2(n15455), .O(n15456) );
  ND2DHD U15719 ( .I1(n15468), .I2(n15456), .O(n15466) );
  AOI22BHD U15720 ( .A1(n7017), .A2(KEY_25), .B1(n13292), .B2(n15457), .O(n15458) );
  OAI112BHD U15721 ( .C1(n10912), .C2(n15460), .A1(n15459), .B1(n15458), .O(n15464) );
  OAI22CHD U15722 ( .A1(n15462), .A2(n15513), .B1(n15512), .B2(n15461), .O(n15463) );
  OAI112BHD U15723 ( .C1(n15468), .C2(n15467), .A1(n15466), .B1(n15465), .O(n6102) );
  AOI22BHD U15724 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _103), .B1(n15504), .B2(_i_CLEFIA128_keyK _39), .O(n15480) );
  AO22CHD U15725 ( .A1(n7045), .A2(n15469), .B1(n15504), .B2(n8626), .O(n15470) );
  AOI22BHD U15726 ( .A1(n7017), .A2(KEY_71), .B1(n13292), .B2(n15471), .O(n15472) );
  OAI112BHD U15727 ( .C1(n10912), .C2(n15474), .A1(n15473), .B1(n15472), .O(n15477) );
  OAI22CHD U15728 ( .A1(n15475), .A2(n15513), .B1(n15512), .B2(n15483), .O(n15476) );
  NR2CHD U15729 ( .I1(n15477), .I2(n15476), .O(n15478) );
  OAI112BHD U15730 ( .C1(n15481), .C2(n15480), .A1(n15479), .B1(n15478), .O(n6151) );
  AOI22BHD U15731 ( .A1(n15492), .A2(DIN_103), .B1(n7017), .B2(KEY_103), .O(n15482) );
  OAI112BHD U15732 ( .C1(n15486), .C2(n11129), .A1(n15485), .B1(n15484), .O(n6197) );
  AOI22BHD U15733 ( .A1(n15492), .A2(DIN_115), .B1(n7017), .B2(KEY_115), .O(n15487) );
  AOI22BHD U15734 ( .A1(n15492), .A2(DIN_51), .B1(n7017), .B2(KEY_51), .O(n15490) );
  AOI22BHD U15735 ( .A1(n15492), .A2(DIN_62), .B1(n7017), .B2(KEY_62), .O(n15493) );
  OAI112BHD U15736 ( .C1(n15503), .C2(n15513), .A1(n15496), .B1(n15495), .O(n6188) );
  AOI22BHD U15737 ( .A1(n15492), .A2(DIN_126), .B1(n7017), .B2(KEY_126), .O(n15497) );
  OAI112BHD U15738 ( .C1(n15503), .C2(n11129), .A1(n15502), .B1(n15501), .O(n6220) );
  AOI22BHD U15739 ( .A1(n7045), .A2(_i_CLEFIA128_keyK _64), .B1(n15504), .B2(_i_CLEFIA128_keyK _0), .O(n15519) );
  AO22CHD U15740 ( .A1(n7045), .A2(n15505), .B1(n15504), .B2(n8777), .O(n15506) );
  AOI22BHD U15741 ( .A1(n7017), .A2(KEY_0), .B1(n13292), .B2(n15507), .O(n15508) );
  OAI112BHD U15742 ( .C1(n10912), .C2(n15510), .A1(n15509), .B1(n15508), .O(n15516) );
  OAI22CHD U15743 ( .A1(n15514), .A2(n15513), .B1(n15512), .B2(n15511), .O(n15515) );
  OAI112BHD U15744 ( .C1(n15520), .C2(n15519), .A1(n15518), .B1(n15517), .O(n6158) );
endmodule
