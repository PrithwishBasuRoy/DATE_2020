module SIMON_enc ( Kin, Din, Dout, Krdy, Drdy, Kvld, Dvld, EN, BSY, CLK, RSTn );
  input [63:0] Kin;
  input [31:0] Din;
  output [31:0] Dout;
  input Krdy, Drdy, EN, CLK, RSTn;
  output Kvld, Dvld, BSY;
  wire   sel, \keyexpantion/N27 , \keyexpantion/N26 , n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857;
  wire   [31:0] rnd;
  wire   [31:0] dat_next;
  wire   [63:0] rkey_next;
  wire   [63:0] rkey;
  wire   [63:0] key;
  assign Dout[31] = dat_next[15];
  assign Dout[30] = dat_next[14];
  assign Dout[29] = dat_next[13];
  assign Dout[28] = dat_next[12];
  assign Dout[27] = dat_next[11];
  assign Dout[26] = dat_next[10];
  assign Dout[25] = dat_next[9];
  assign Dout[24] = dat_next[8];
  assign Dout[23] = dat_next[7];
  assign Dout[22] = dat_next[6];
  assign Dout[21] = dat_next[5];
  assign Dout[20] = dat_next[4];
  assign Dout[19] = dat_next[3];
  assign Dout[18] = dat_next[2];
  assign Dout[17] = dat_next[1];
  assign Dout[16] = dat_next[0];

  QDFFRBHHD Kvld_reg ( .D(n483), .CK(CLK), .RB(RSTn), .Q(Kvld) );
  QDFFRBHHD sel_reg ( .D(n482), .CK(CLK), .RB(RSTn), .Q(sel) );
  QDFFRBHHD Dvld_reg ( .D(n481), .CK(CLK), .RB(RSTn), .Q(Dvld) );
  QDFFRBHHD BSY_reg ( .D(n480), .CK(CLK), .RB(RSTn), .Q(BSY) );
  QDFFRBHHD \rkey_reg[0]  ( .D(n479), .CK(CLK), .RB(RSTn), .Q(rkey[0]) );
  QDFFRBHHD \rkey_reg[48]  ( .D(n478), .CK(CLK), .RB(RSTn), .Q(rkey_next[32])
         );
  QDFFRBHHD \rkey_reg[32]  ( .D(n477), .CK(CLK), .RB(RSTn), .Q(rkey_next[16])
         );
  QDFFRBHHD \rkey_reg[16]  ( .D(n476), .CK(CLK), .RB(RSTn), .Q(rkey_next[0])
         );
  QDFFRBHHD \rkey_reg[61]  ( .D(n475), .CK(CLK), .RB(RSTn), .Q(rkey_next[45])
         );
  QDFFRBHHD \rkey_reg[45]  ( .D(n474), .CK(CLK), .RB(RSTn), .Q(rkey_next[29])
         );
  QDFFRBHHD \rkey_reg[29]  ( .D(n473), .CK(CLK), .RB(RSTn), .Q(rkey_next[13])
         );
  QDFFRBHHD \rkey_reg[13]  ( .D(n472), .CK(CLK), .RB(RSTn), .Q(rkey[13]) );
  QDFFRBHHD \rkey_reg[58]  ( .D(n471), .CK(CLK), .RB(RSTn), .Q(rkey_next[42])
         );
  QDFFRBHHD \rkey_reg[42]  ( .D(n470), .CK(CLK), .RB(RSTn), .Q(rkey_next[26])
         );
  QDFFRBHHD \rkey_reg[26]  ( .D(n469), .CK(CLK), .RB(RSTn), .Q(rkey_next[10])
         );
  QDFFRBHHD \rkey_reg[10]  ( .D(n468), .CK(CLK), .RB(RSTn), .Q(rkey[10]) );
  QDFFRBHHD \rkey_reg[55]  ( .D(n467), .CK(CLK), .RB(RSTn), .Q(rkey_next[39])
         );
  QDFFRBHHD \rkey_reg[39]  ( .D(n466), .CK(CLK), .RB(RSTn), .Q(rkey_next[23])
         );
  QDFFRBHHD \rkey_reg[23]  ( .D(n465), .CK(CLK), .RB(RSTn), .Q(rkey_next[7])
         );
  QDFFRBHHD \rkey_reg[7]  ( .D(n464), .CK(CLK), .RB(RSTn), .Q(rkey[7]) );
  QDFFRBHHD \rkey_reg[52]  ( .D(n463), .CK(CLK), .RB(RSTn), .Q(rkey_next[36])
         );
  QDFFRBHHD \rkey_reg[36]  ( .D(n462), .CK(CLK), .RB(RSTn), .Q(rkey_next[20])
         );
  QDFFRBHHD \rkey_reg[20]  ( .D(n461), .CK(CLK), .RB(RSTn), .Q(rkey_next[4])
         );
  QDFFRBHHD \rkey_reg[4]  ( .D(n460), .CK(CLK), .RB(RSTn), .Q(rkey[4]) );
  QDFFRBHHD \rkey_reg[49]  ( .D(n459), .CK(CLK), .RB(RSTn), .Q(rkey_next[33])
         );
  QDFFRBHHD \rkey_reg[33]  ( .D(n458), .CK(CLK), .RB(RSTn), .Q(rkey_next[17])
         );
  QDFFRBHHD \rkey_reg[17]  ( .D(n457), .CK(CLK), .RB(RSTn), .Q(rkey_next[1])
         );
  QDFFRBHHD \rkey_reg[1]  ( .D(n456), .CK(CLK), .RB(RSTn), .Q(rkey[1]) );
  QDFFRBHHD \rkey_reg[62]  ( .D(n455), .CK(CLK), .RB(RSTn), .Q(rkey_next[46])
         );
  QDFFRBHHD \rkey_reg[46]  ( .D(n454), .CK(CLK), .RB(RSTn), .Q(rkey_next[30])
         );
  QDFFRBHHD \rkey_reg[30]  ( .D(n453), .CK(CLK), .RB(RSTn), .Q(rkey_next[14])
         );
  QDFFRBHHD \rkey_reg[14]  ( .D(n452), .CK(CLK), .RB(RSTn), .Q(rkey[14]) );
  QDFFRBHHD \rkey_reg[59]  ( .D(n451), .CK(CLK), .RB(RSTn), .Q(rkey_next[43])
         );
  QDFFRBHHD \rkey_reg[43]  ( .D(n450), .CK(CLK), .RB(RSTn), .Q(rkey_next[27])
         );
  QDFFRBHHD \rkey_reg[27]  ( .D(n449), .CK(CLK), .RB(RSTn), .Q(rkey_next[11])
         );
  QDFFRBHHD \rkey_reg[11]  ( .D(n448), .CK(CLK), .RB(RSTn), .Q(rkey[11]) );
  QDFFRBHHD \rkey_reg[56]  ( .D(n447), .CK(CLK), .RB(RSTn), .Q(rkey_next[40])
         );
  QDFFRBHHD \rkey_reg[40]  ( .D(n446), .CK(CLK), .RB(RSTn), .Q(rkey_next[24])
         );
  QDFFRBHHD \rkey_reg[24]  ( .D(n445), .CK(CLK), .RB(RSTn), .Q(rkey_next[8])
         );
  QDFFRBHHD \rkey_reg[8]  ( .D(n444), .CK(CLK), .RB(RSTn), .Q(rkey[8]) );
  QDFFRBHHD \rkey_reg[53]  ( .D(n443), .CK(CLK), .RB(RSTn), .Q(rkey_next[37])
         );
  QDFFRBHHD \rkey_reg[37]  ( .D(n442), .CK(CLK), .RB(RSTn), .Q(rkey_next[21])
         );
  QDFFRBHHD \rkey_reg[21]  ( .D(n441), .CK(CLK), .RB(RSTn), .Q(rkey_next[5])
         );
  QDFFRBHHD \rkey_reg[5]  ( .D(n440), .CK(CLK), .RB(RSTn), .Q(rkey[5]) );
  QDFFRBHHD \rkey_reg[50]  ( .D(n439), .CK(CLK), .RB(RSTn), .Q(rkey_next[34])
         );
  QDFFRBHHD \rkey_reg[34]  ( .D(n438), .CK(CLK), .RB(RSTn), .Q(rkey_next[18])
         );
  QDFFRBHHD \rkey_reg[18]  ( .D(n437), .CK(CLK), .RB(RSTn), .Q(rkey_next[2])
         );
  QDFFRBHHD \rkey_reg[2]  ( .D(n436), .CK(CLK), .RB(RSTn), .Q(rkey[2]) );
  QDFFRBHHD \rkey_reg[63]  ( .D(n435), .CK(CLK), .RB(RSTn), .Q(rkey_next[47])
         );
  QDFFRBHHD \rkey_reg[47]  ( .D(n434), .CK(CLK), .RB(RSTn), .Q(rkey_next[31])
         );
  QDFFRBHHD \rkey_reg[31]  ( .D(n433), .CK(CLK), .RB(RSTn), .Q(rkey_next[15])
         );
  QDFFRBHHD \rkey_reg[15]  ( .D(n432), .CK(CLK), .RB(RSTn), .Q(rkey[15]) );
  QDFFRBHHD \rkey_reg[60]  ( .D(n431), .CK(CLK), .RB(RSTn), .Q(rkey_next[44])
         );
  QDFFRBHHD \rkey_reg[44]  ( .D(n430), .CK(CLK), .RB(RSTn), .Q(rkey_next[28])
         );
  QDFFRBHHD \rkey_reg[28]  ( .D(n429), .CK(CLK), .RB(RSTn), .Q(rkey_next[12])
         );
  QDFFRBHHD \rkey_reg[12]  ( .D(n428), .CK(CLK), .RB(RSTn), .Q(rkey[12]) );
  QDFFRBHHD \rkey_reg[57]  ( .D(n427), .CK(CLK), .RB(RSTn), .Q(rkey_next[41])
         );
  QDFFRBHHD \rkey_reg[41]  ( .D(n426), .CK(CLK), .RB(RSTn), .Q(rkey_next[25])
         );
  QDFFRBHHD \rkey_reg[25]  ( .D(n425), .CK(CLK), .RB(RSTn), .Q(rkey_next[9])
         );
  QDFFRBHHD \rkey_reg[9]  ( .D(n424), .CK(CLK), .RB(RSTn), .Q(rkey[9]) );
  QDFFRBHHD \rkey_reg[54]  ( .D(n423), .CK(CLK), .RB(RSTn), .Q(rkey_next[38])
         );
  QDFFRBHHD \rkey_reg[38]  ( .D(n422), .CK(CLK), .RB(RSTn), .Q(rkey_next[22])
         );
  QDFFRBHHD \rkey_reg[22]  ( .D(n421), .CK(CLK), .RB(RSTn), .Q(rkey_next[6])
         );
  QDFFRBHHD \rkey_reg[6]  ( .D(n420), .CK(CLK), .RB(RSTn), .Q(rkey[6]) );
  QDFFRBHHD \rkey_reg[51]  ( .D(n419), .CK(CLK), .RB(RSTn), .Q(rkey_next[35])
         );
  QDFFRBHHD \rkey_reg[35]  ( .D(n418), .CK(CLK), .RB(RSTn), .Q(rkey_next[19])
         );
  QDFFRBHHD \rkey_reg[19]  ( .D(n417), .CK(CLK), .RB(RSTn), .Q(rkey_next[3])
         );
  QDFFRBHHD \rkey_reg[3]  ( .D(n416), .CK(CLK), .RB(RSTn), .Q(rkey[3]) );
  QDFFRBHHD \rnd_reg[1]  ( .D(n610), .CK(CLK), .RB(RSTn), .Q(
        \keyexpantion/N27 ) );
  QDFFRBHHD \rnd_reg[2]  ( .D(n609), .CK(CLK), .RB(RSTn), .Q(rnd[2]) );
  QDFFRBHHD \rnd_reg[3]  ( .D(n608), .CK(CLK), .RB(RSTn), .Q(rnd[3]) );
  QDFFRBHHD \rnd_reg[4]  ( .D(n607), .CK(CLK), .RB(RSTn), .Q(rnd[4]) );
  QDFFRBHHD \rnd_reg[5]  ( .D(n606), .CK(CLK), .RB(RSTn), .Q(rnd[5]) );
  QDFFRBHHD \rnd_reg[6]  ( .D(n605), .CK(CLK), .RB(RSTn), .Q(rnd[6]) );
  QDFFRBHHD \rnd_reg[7]  ( .D(n604), .CK(CLK), .RB(RSTn), .Q(rnd[7]) );
  QDFFRBHHD \rnd_reg[8]  ( .D(n603), .CK(CLK), .RB(RSTn), .Q(rnd[8]) );
  QDFFRBHHD \rnd_reg[9]  ( .D(n602), .CK(CLK), .RB(RSTn), .Q(rnd[9]) );
  QDFFRBHHD \rnd_reg[10]  ( .D(n601), .CK(CLK), .RB(RSTn), .Q(rnd[10]) );
  QDFFRBHHD \rnd_reg[11]  ( .D(n600), .CK(CLK), .RB(RSTn), .Q(rnd[11]) );
  QDFFRBHHD \rnd_reg[12]  ( .D(n599), .CK(CLK), .RB(RSTn), .Q(rnd[12]) );
  QDFFRBHHD \rnd_reg[13]  ( .D(n598), .CK(CLK), .RB(RSTn), .Q(rnd[13]) );
  QDFFRBHHD \rnd_reg[14]  ( .D(n597), .CK(CLK), .RB(RSTn), .Q(rnd[14]) );
  QDFFRBHHD \rnd_reg[15]  ( .D(n596), .CK(CLK), .RB(RSTn), .Q(rnd[15]) );
  QDFFRBHHD \rnd_reg[16]  ( .D(n595), .CK(CLK), .RB(RSTn), .Q(rnd[16]) );
  QDFFRBHHD \rnd_reg[17]  ( .D(n594), .CK(CLK), .RB(RSTn), .Q(rnd[17]) );
  QDFFRBHHD \rnd_reg[18]  ( .D(n593), .CK(CLK), .RB(RSTn), .Q(rnd[18]) );
  QDFFRBHHD \rnd_reg[19]  ( .D(n592), .CK(CLK), .RB(RSTn), .Q(rnd[19]) );
  QDFFRBHHD \rnd_reg[20]  ( .D(n591), .CK(CLK), .RB(RSTn), .Q(rnd[20]) );
  QDFFRBHHD \rnd_reg[21]  ( .D(n590), .CK(CLK), .RB(RSTn), .Q(rnd[21]) );
  QDFFRBHHD \rnd_reg[22]  ( .D(n589), .CK(CLK), .RB(RSTn), .Q(rnd[22]) );
  QDFFRBHHD \rnd_reg[23]  ( .D(n588), .CK(CLK), .RB(RSTn), .Q(rnd[23]) );
  QDFFRBHHD \rnd_reg[24]  ( .D(n587), .CK(CLK), .RB(RSTn), .Q(rnd[24]) );
  QDFFRBHHD \rnd_reg[25]  ( .D(n586), .CK(CLK), .RB(RSTn), .Q(rnd[25]) );
  QDFFRBHHD \rnd_reg[26]  ( .D(n585), .CK(CLK), .RB(RSTn), .Q(rnd[26]) );
  QDFFRBHHD \rnd_reg[27]  ( .D(n584), .CK(CLK), .RB(RSTn), .Q(rnd[27]) );
  QDFFRBHHD \rnd_reg[28]  ( .D(n583), .CK(CLK), .RB(RSTn), .Q(rnd[28]) );
  QDFFRBHHD \rnd_reg[29]  ( .D(n582), .CK(CLK), .RB(RSTn), .Q(rnd[29]) );
  QDFFRBHHD \rnd_reg[30]  ( .D(n581), .CK(CLK), .RB(RSTn), .Q(rnd[30]) );
  QDFFRBHHD \rnd_reg[31]  ( .D(n612), .CK(CLK), .RB(RSTn), .Q(rnd[31]) );
  QDFFRBHHD \key_reg[63]  ( .D(n580), .CK(CLK), .RB(RSTn), .Q(key[63]) );
  QDFFRBHHD \key_reg[62]  ( .D(n579), .CK(CLK), .RB(RSTn), .Q(key[62]) );
  QDFFRBHHD \key_reg[61]  ( .D(n578), .CK(CLK), .RB(RSTn), .Q(key[61]) );
  QDFFRBHHD \key_reg[60]  ( .D(n577), .CK(CLK), .RB(RSTn), .Q(key[60]) );
  QDFFRBHHD \key_reg[59]  ( .D(n576), .CK(CLK), .RB(RSTn), .Q(key[59]) );
  QDFFRBHHD \key_reg[58]  ( .D(n575), .CK(CLK), .RB(RSTn), .Q(key[58]) );
  QDFFRBHHD \key_reg[57]  ( .D(n574), .CK(CLK), .RB(RSTn), .Q(key[57]) );
  QDFFRBHHD \key_reg[56]  ( .D(n573), .CK(CLK), .RB(RSTn), .Q(key[56]) );
  QDFFRBHHD \key_reg[55]  ( .D(n572), .CK(CLK), .RB(RSTn), .Q(key[55]) );
  QDFFRBHHD \key_reg[54]  ( .D(n571), .CK(CLK), .RB(RSTn), .Q(key[54]) );
  QDFFRBHHD \key_reg[53]  ( .D(n570), .CK(CLK), .RB(RSTn), .Q(key[53]) );
  QDFFRBHHD \key_reg[52]  ( .D(n569), .CK(CLK), .RB(RSTn), .Q(key[52]) );
  QDFFRBHHD \key_reg[51]  ( .D(n568), .CK(CLK), .RB(RSTn), .Q(key[51]) );
  QDFFRBHHD \key_reg[50]  ( .D(n567), .CK(CLK), .RB(RSTn), .Q(key[50]) );
  QDFFRBHHD \key_reg[49]  ( .D(n566), .CK(CLK), .RB(RSTn), .Q(key[49]) );
  QDFFRBHHD \key_reg[48]  ( .D(n565), .CK(CLK), .RB(RSTn), .Q(key[48]) );
  QDFFRBHHD \key_reg[47]  ( .D(n564), .CK(CLK), .RB(RSTn), .Q(key[47]) );
  QDFFRBHHD \key_reg[46]  ( .D(n563), .CK(CLK), .RB(RSTn), .Q(key[46]) );
  QDFFRBHHD \key_reg[45]  ( .D(n562), .CK(CLK), .RB(RSTn), .Q(key[45]) );
  QDFFRBHHD \key_reg[44]  ( .D(n561), .CK(CLK), .RB(RSTn), .Q(key[44]) );
  QDFFRBHHD \key_reg[43]  ( .D(n560), .CK(CLK), .RB(RSTn), .Q(key[43]) );
  QDFFRBHHD \key_reg[42]  ( .D(n559), .CK(CLK), .RB(RSTn), .Q(key[42]) );
  QDFFRBHHD \key_reg[41]  ( .D(n558), .CK(CLK), .RB(RSTn), .Q(key[41]) );
  QDFFRBHHD \key_reg[40]  ( .D(n557), .CK(CLK), .RB(RSTn), .Q(key[40]) );
  QDFFRBHHD \key_reg[39]  ( .D(n556), .CK(CLK), .RB(RSTn), .Q(key[39]) );
  QDFFRBHHD \key_reg[38]  ( .D(n555), .CK(CLK), .RB(RSTn), .Q(key[38]) );
  QDFFRBHHD \key_reg[37]  ( .D(n554), .CK(CLK), .RB(RSTn), .Q(key[37]) );
  QDFFRBHHD \key_reg[36]  ( .D(n553), .CK(CLK), .RB(RSTn), .Q(key[36]) );
  QDFFRBHHD \key_reg[35]  ( .D(n552), .CK(CLK), .RB(RSTn), .Q(key[35]) );
  QDFFRBHHD \key_reg[34]  ( .D(n551), .CK(CLK), .RB(RSTn), .Q(key[34]) );
  QDFFRBHHD \key_reg[33]  ( .D(n550), .CK(CLK), .RB(RSTn), .Q(key[33]) );
  QDFFRBHHD \key_reg[32]  ( .D(n549), .CK(CLK), .RB(RSTn), .Q(key[32]) );
  QDFFRBHHD \key_reg[31]  ( .D(n548), .CK(CLK), .RB(RSTn), .Q(key[31]) );
  QDFFRBHHD \key_reg[30]  ( .D(n547), .CK(CLK), .RB(RSTn), .Q(key[30]) );
  QDFFRBHHD \key_reg[29]  ( .D(n546), .CK(CLK), .RB(RSTn), .Q(key[29]) );
  QDFFRBHHD \key_reg[28]  ( .D(n545), .CK(CLK), .RB(RSTn), .Q(key[28]) );
  QDFFRBHHD \key_reg[27]  ( .D(n544), .CK(CLK), .RB(RSTn), .Q(key[27]) );
  QDFFRBHHD \key_reg[26]  ( .D(n543), .CK(CLK), .RB(RSTn), .Q(key[26]) );
  QDFFRBHHD \key_reg[25]  ( .D(n542), .CK(CLK), .RB(RSTn), .Q(key[25]) );
  QDFFRBHHD \key_reg[24]  ( .D(n541), .CK(CLK), .RB(RSTn), .Q(key[24]) );
  QDFFRBHHD \key_reg[23]  ( .D(n540), .CK(CLK), .RB(RSTn), .Q(key[23]) );
  QDFFRBHHD \key_reg[22]  ( .D(n539), .CK(CLK), .RB(RSTn), .Q(key[22]) );
  QDFFRBHHD \key_reg[21]  ( .D(n538), .CK(CLK), .RB(RSTn), .Q(key[21]) );
  QDFFRBHHD \key_reg[20]  ( .D(n537), .CK(CLK), .RB(RSTn), .Q(key[20]) );
  QDFFRBHHD \key_reg[19]  ( .D(n536), .CK(CLK), .RB(RSTn), .Q(key[19]) );
  QDFFRBHHD \key_reg[18]  ( .D(n535), .CK(CLK), .RB(RSTn), .Q(key[18]) );
  QDFFRBHHD \key_reg[17]  ( .D(n534), .CK(CLK), .RB(RSTn), .Q(key[17]) );
  QDFFRBHHD \key_reg[16]  ( .D(n533), .CK(CLK), .RB(RSTn), .Q(key[16]) );
  QDFFRBHHD \key_reg[15]  ( .D(n532), .CK(CLK), .RB(RSTn), .Q(key[15]) );
  QDFFRBHHD \key_reg[14]  ( .D(n531), .CK(CLK), .RB(RSTn), .Q(key[14]) );
  QDFFRBHHD \key_reg[13]  ( .D(n530), .CK(CLK), .RB(RSTn), .Q(key[13]) );
  QDFFRBHHD \key_reg[12]  ( .D(n529), .CK(CLK), .RB(RSTn), .Q(key[12]) );
  QDFFRBHHD \key_reg[11]  ( .D(n528), .CK(CLK), .RB(RSTn), .Q(key[11]) );
  QDFFRBHHD \key_reg[10]  ( .D(n527), .CK(CLK), .RB(RSTn), .Q(key[10]) );
  QDFFRBHHD \key_reg[9]  ( .D(n526), .CK(CLK), .RB(RSTn), .Q(key[9]) );
  QDFFRBHHD \key_reg[8]  ( .D(n525), .CK(CLK), .RB(RSTn), .Q(key[8]) );
  QDFFRBHHD \key_reg[7]  ( .D(n524), .CK(CLK), .RB(RSTn), .Q(key[7]) );
  QDFFRBHHD \key_reg[6]  ( .D(n523), .CK(CLK), .RB(RSTn), .Q(key[6]) );
  QDFFRBHHD \key_reg[5]  ( .D(n522), .CK(CLK), .RB(RSTn), .Q(key[5]) );
  QDFFRBHHD \key_reg[4]  ( .D(n521), .CK(CLK), .RB(RSTn), .Q(key[4]) );
  QDFFRBHHD \key_reg[3]  ( .D(n520), .CK(CLK), .RB(RSTn), .Q(key[3]) );
  QDFFRBHHD \key_reg[2]  ( .D(n519), .CK(CLK), .RB(RSTn), .Q(key[2]) );
  QDFFRBHHD \key_reg[1]  ( .D(n518), .CK(CLK), .RB(RSTn), .Q(key[1]) );
  QDFFRBHHD \key_reg[0]  ( .D(n517), .CK(CLK), .RB(RSTn), .Q(key[0]) );
  QDFFRBHHD \dat_reg[16]  ( .D(n500), .CK(CLK), .RB(RSTn), .Q(dat_next[0]) );
  QDFFRBHHD \dat_reg[0]  ( .D(n516), .CK(CLK), .RB(RSTn), .Q(Dout[0]) );
  QDFFRBHHD \dat_reg[24]  ( .D(n492), .CK(CLK), .RB(RSTn), .Q(dat_next[8]) );
  QDFFRBHHD \dat_reg[8]  ( .D(n508), .CK(CLK), .RB(RSTn), .Q(Dout[8]) );
  QDFFRBHHD \dat_reg[26]  ( .D(n490), .CK(CLK), .RB(RSTn), .Q(dat_next[10]) );
  QDFFRBHHD \dat_reg[10]  ( .D(n506), .CK(CLK), .RB(RSTn), .Q(Dout[10]) );
  QDFFRBHHD \dat_reg[28]  ( .D(n488), .CK(CLK), .RB(RSTn), .Q(dat_next[12]) );
  QDFFRBHHD \dat_reg[12]  ( .D(n504), .CK(CLK), .RB(RSTn), .Q(Dout[12]) );
  QDFFRBHHD \dat_reg[30]  ( .D(n486), .CK(CLK), .RB(RSTn), .Q(dat_next[14]) );
  QDFFRBHHD \dat_reg[14]  ( .D(n502), .CK(CLK), .RB(RSTn), .Q(Dout[14]) );
  QDFFRBHHD \dat_reg[31]  ( .D(n484), .CK(CLK), .RB(RSTn), .Q(dat_next[15]) );
  QDFFRBHHD \dat_reg[15]  ( .D(n501), .CK(CLK), .RB(RSTn), .Q(Dout[15]) );
  QDFFRBHHD \dat_reg[23]  ( .D(n493), .CK(CLK), .RB(RSTn), .Q(dat_next[7]) );
  QDFFRBHHD \dat_reg[7]  ( .D(n509), .CK(CLK), .RB(RSTn), .Q(Dout[7]) );
  QDFFRBHHD \dat_reg[25]  ( .D(n491), .CK(CLK), .RB(RSTn), .Q(dat_next[9]) );
  QDFFRBHHD \dat_reg[9]  ( .D(n507), .CK(CLK), .RB(RSTn), .Q(Dout[9]) );
  QDFFRBHHD \dat_reg[17]  ( .D(n499), .CK(CLK), .RB(RSTn), .Q(dat_next[1]) );
  QDFFRBHHD \dat_reg[1]  ( .D(n515), .CK(CLK), .RB(RSTn), .Q(Dout[1]) );
  QDFFRBHHD \dat_reg[18]  ( .D(n498), .CK(CLK), .RB(RSTn), .Q(dat_next[2]) );
  QDFFRBHHD \dat_reg[2]  ( .D(n514), .CK(CLK), .RB(RSTn), .Q(Dout[2]) );
  QDFFRBHHD \dat_reg[27]  ( .D(n489), .CK(CLK), .RB(RSTn), .Q(dat_next[11]) );
  QDFFRBHHD \dat_reg[11]  ( .D(n505), .CK(CLK), .RB(RSTn), .Q(Dout[11]) );
  QDFFRBHHD \dat_reg[19]  ( .D(n497), .CK(CLK), .RB(RSTn), .Q(dat_next[3]) );
  QDFFRBHHD \dat_reg[3]  ( .D(n513), .CK(CLK), .RB(RSTn), .Q(Dout[3]) );
  QDFFRBHHD \dat_reg[20]  ( .D(n496), .CK(CLK), .RB(RSTn), .Q(dat_next[4]) );
  QDFFRBHHD \dat_reg[4]  ( .D(n512), .CK(CLK), .RB(RSTn), .Q(Dout[4]) );
  QDFFRBHHD \dat_reg[29]  ( .D(n487), .CK(CLK), .RB(RSTn), .Q(dat_next[13]) );
  QDFFRBHHD \dat_reg[13]  ( .D(n503), .CK(CLK), .RB(RSTn), .Q(Dout[13]) );
  QDFFRBHHD \dat_reg[21]  ( .D(n495), .CK(CLK), .RB(RSTn), .Q(dat_next[5]) );
  QDFFRBHHD \dat_reg[5]  ( .D(n511), .CK(CLK), .RB(RSTn), .Q(Dout[5]) );
  QDFFRBHHD \dat_reg[22]  ( .D(n494), .CK(CLK), .RB(RSTn), .Q(dat_next[6]) );
  QDFFRBHHD \dat_reg[6]  ( .D(n510), .CK(CLK), .RB(RSTn), .Q(Dout[6]) );
  DFFSBEHD \rnd_reg[0]  ( .D(n611), .CK(CLK), .SB(RSTn), .Q(\keyexpantion/N26 ), .QB(n1857) );
  INVDHD U616 ( .I(EN), .O(n1584) );
  INVDHD U617 ( .I(n734), .O(n652) );
  NR2EHD U618 ( .I1(n735), .I2(n724), .O(n723) );
  INVDHD U619 ( .I(n1291), .O(n1289) );
  XNR2EHD U620 ( .I1(n1217), .I2(n1216), .O(n1236) );
  INVDHD U621 ( .I(n1021), .O(n1028) );
  XNR2EHD U622 ( .I1(n1098), .I2(n1100), .O(n627) );
  INVDHD U623 ( .I(n681), .O(n849) );
  INVDHD U624 ( .I(n1250), .O(n660) );
  XNR2HHD U625 ( .I1(n1069), .I2(n1202), .O(n1118) );
  ND2CHD U626 ( .I1(n1006), .I2(rnd[28]), .O(n1009) );
  XOR2EHD U627 ( .I1(rnd[25]), .I2(n1073), .O(n1072) );
  INVGHD U628 ( .I(n1005), .O(n1092) );
  XNR2HHD U629 ( .I1(n1091), .I2(n1005), .O(n1144) );
  NR2GHD U630 ( .I1(n987), .I2(n1062), .O(n1000) );
  INVHHD U631 ( .I(n898), .O(n1061) );
  INVDHD U632 ( .I(n982), .O(n755) );
  XNR2HHD U633 ( .I1(rnd[15]), .I2(n694), .O(n1039) );
  ND2DHD U634 ( .I1(n749), .I2(n787), .O(n748) );
  INVGHD U635 ( .I(rnd[2]), .O(n1579) );
  BUFCKIHD U636 ( .I(n975), .O(n632) );
  INVGHD U637 ( .I(rnd[19]), .O(n1561) );
  INVGHD U638 ( .I(rnd[20]), .O(n1562) );
  INVLHD U639 ( .I(rnd[14]), .O(n1350) );
  XNR2EHD U640 ( .I1(n1108), .I2(n621), .O(n1132) );
  ND2HHD U641 ( .I1(n750), .I2(n748), .O(n1140) );
  XNR2HHD U642 ( .I1(rnd[29]), .I2(n1113), .O(n1252) );
  BUFEHD U643 ( .I(n1330), .O(n1852) );
  ND2DHD U644 ( .I1(n1349), .I2(EN), .O(n1570) );
  INVKHD U645 ( .I(n868), .O(n917) );
  INVLHD U646 ( .I(n1034), .O(n768) );
  ND2HHD U647 ( .I1(n1201), .I2(n1200), .O(n1235) );
  ND2HHD U648 ( .I1(n1255), .I2(n1114), .O(n1065) );
  INVDHD U649 ( .I(n1150), .O(n1153) );
  NR2GHD U650 ( .I1(rnd[19]), .I2(rnd[18]), .O(n934) );
  NR2EHD U651 ( .I1(n1148), .I2(n780), .O(n779) );
  MAO222EHD U652 ( .A1(n1147), .B1(n1146), .C1(n1145), .O(n1148) );
  NR2BHD U653 ( .I1(n789), .I2(n869), .O(n786) );
  ND2HHD U654 ( .I1(n1104), .I2(n1103), .O(n1151) );
  INVCHD U655 ( .I(n1047), .O(n1048) );
  AN2HHD U656 ( .I1(n1074), .I2(n719), .O(n1047) );
  INVGHD U657 ( .I(n758), .O(n733) );
  ND2DHD U658 ( .I1(n1030), .I2(n1031), .O(n741) );
  INVCKGHD U659 ( .I(n632), .O(n1319) );
  INVCKGHD U660 ( .I(n1222), .O(n683) );
  ND2HHD U661 ( .I1(n904), .I2(n923), .O(n907) );
  NR2CHD U662 ( .I1(n918), .I2(n1315), .O(n919) );
  OA12EHD U663 ( .B1(n992), .B2(n996), .A1(n995), .O(n1111) );
  XNR2KHD U664 ( .I1(n1082), .I2(n1081), .O(n1087) );
  ND2HHD U665 ( .I1(n892), .I2(n891), .O(n906) );
  INVGHD U666 ( .I(n1163), .O(n614) );
  AOI22BHD U667 ( .A1(Din[16]), .A2(n1573), .B1(n1571), .B2(dat_next[0]), .O(
        n1299) );
  ND2DHD U668 ( .I1(n1298), .I2(EN), .O(n1571) );
  NR2CHD U669 ( .I1(n1577), .I2(n1578), .O(n1845) );
  NR2CHD U670 ( .I1(n1579), .I2(n1578), .O(n1851) );
  MXL2CHD U671 ( .A(n1561), .B(n1562), .S(n1570), .OB(n591) );
  MXL2CHD U672 ( .A(n1560), .B(n1561), .S(n1570), .OB(n592) );
  XNR2CHD U673 ( .I1(rnd[7]), .I2(n746), .O(n745) );
  AN2HHD U674 ( .I1(n1297), .I2(n1295), .O(n1572) );
  ND2DHD U675 ( .I1(n1583), .I2(n1553), .O(n1578) );
  AN2EHD U676 ( .I1(\keyexpantion/N27 ), .I2(n1583), .O(n1844) );
  ND2DHD U677 ( .I1(n1294), .I2(\keyexpantion/N26 ), .O(n1297) );
  NR2CHD U678 ( .I1(n1328), .I2(\keyexpantion/N26 ), .O(n1583) );
  INVDHD U679 ( .I(\keyexpantion/N27 ), .O(n1553) );
  ND2DHD U680 ( .I1(\keyexpantion/N26 ), .I2(n1348), .O(n1349) );
  INVGHD U681 ( .I(rnd[6]), .O(n914) );
  NR2CHD U682 ( .I1(Drdy), .I2(n1584), .O(n1295) );
  ND2DHD U683 ( .I1(n1327), .I2(EN), .O(n1328) );
  AN2EHD U684 ( .I1(EN), .I2(Drdy), .O(n1573) );
  AN2HHD U685 ( .I1(EN), .I2(Krdy), .O(n1807) );
  XNR2HHD U686 ( .I1(n1129), .I2(n1126), .O(n780) );
  OR2EHD U687 ( .I1(n1022), .I2(n785), .O(n617) );
  ND2HHD U688 ( .I1(n861), .I2(n860), .O(n862) );
  BUFLHD U689 ( .I(n975), .O(n878) );
  ND2HHD U690 ( .I1(n740), .I2(n991), .O(n998) );
  ND2HHD U691 ( .I1(n1115), .I2(n1202), .O(n848) );
  NR2IHD U692 ( .I1(rnd[14]), .I2(n1115), .O(n681) );
  INVGHD U693 ( .I(n1115), .O(n1255) );
  INVCKGHD U694 ( .I(n965), .O(n966) );
  XNR2KHD U695 ( .I1(rnd[31]), .I2(n876), .O(n896) );
  NR2GHD U696 ( .I1(\keyexpantion/N26 ), .I2(n1137), .O(n990) );
  INVGHD U697 ( .I(n1143), .O(n997) );
  INVCKGHD U698 ( .I(n1110), .O(n984) );
  NR2CHD U699 ( .I1(n1163), .I2(n758), .O(n757) );
  INVHHD U700 ( .I(n988), .O(n999) );
  INVHHD U701 ( .I(n842), .O(n1329) );
  NR2GHD U702 ( .I1(n852), .I2(n1034), .O(n877) );
  NR2GHD U703 ( .I1(n1033), .I2(n1034), .O(n821) );
  NR2GHD U704 ( .I1(rnd[18]), .I2(n1034), .O(n794) );
  ND2HHD U705 ( .I1(n638), .I2(n637), .O(n959) );
  ND2DHD U706 ( .I1(n882), .I2(n881), .O(n886) );
  INVGHD U707 ( .I(n1114), .O(n1066) );
  NR2EHD U708 ( .I1(n875), .I2(n1034), .O(n876) );
  INVLHD U709 ( .I(n820), .O(n1034) );
  ND2DHD U710 ( .I1(n951), .I2(n997), .O(n955) );
  XNR2HHD U711 ( .I1(n1143), .I2(n698), .O(n1041) );
  NR2EHD U712 ( .I1(n910), .I2(n1034), .O(n773) );
  XNR2HHD U713 ( .I1(n1560), .I2(n1034), .O(n1005) );
  INVDHD U714 ( .I(n1270), .O(n1275) );
  AN2HHD U715 ( .I1(n1272), .I2(n1270), .O(n615) );
  ND2HHD U716 ( .I1(n658), .I2(n1183), .O(n642) );
  ND2DHD U717 ( .I1(n1239), .I2(n1566), .O(n861) );
  INVDHD U718 ( .I(n1215), .O(n1239) );
  ND3CHD U719 ( .I1(n766), .I2(n764), .I3(n765), .O(n763) );
  INVCKGHD U720 ( .I(n765), .O(n762) );
  INVCKGHD U721 ( .I(n879), .O(n856) );
  ND2HHD U722 ( .I1(n739), .I2(n989), .O(n1001) );
  XNR2HHD U723 ( .I1(n1565), .I2(n821), .O(n989) );
  XNR2KHD U724 ( .I1(n1004), .I2(n1003), .O(n1056) );
  XNR2EHD U725 ( .I1(n1064), .I2(n1063), .O(n1082) );
  INVCHD U726 ( .I(n1062), .O(n1063) );
  ND2HHD U727 ( .I1(n751), .I2(n788), .O(n750) );
  ND3CHD U728 ( .I1(n1050), .I2(n1049), .I3(n1048), .O(n1053) );
  XNR2HHD U729 ( .I1(rnd[25]), .I2(n877), .O(n1242) );
  NR2EHD U730 ( .I1(n939), .I2(n938), .O(n940) );
  ND2HHD U731 ( .I1(n701), .I2(n700), .O(n1081) );
  ND2HHD U732 ( .I1(n768), .I2(n1015), .O(n1113) );
  NR2IHD U733 ( .I1(n1061), .I2(n896), .O(n988) );
  NR2EHD U734 ( .I1(rnd[25]), .I2(rnd[24]), .O(n871) );
  ND3CHD U735 ( .I1(n1306), .I2(n865), .I3(n914), .O(n866) );
  NR2GHD U736 ( .I1(n1167), .I2(n668), .O(n667) );
  ND2DHD U737 ( .I1(n1097), .I2(n1096), .O(n742) );
  ND2DHD U738 ( .I1(n1117), .I2(n1118), .O(n1096) );
  ND2KHD U739 ( .I1(n1306), .I2(n943), .O(n932) );
  ND2DHD U740 ( .I1(n1099), .I2(n1072), .O(n700) );
  INVGHD U741 ( .I(n1140), .O(n991) );
  ND2HHD U742 ( .I1(n889), .I2(n888), .O(n892) );
  ND2HHD U743 ( .I1(n1115), .I2(n1066), .O(n1067) );
  AN3EHD U744 ( .I1(n1305), .I2(n1306), .I3(n1561), .O(n832) );
  NR2GHD U745 ( .I1(rnd[17]), .I2(rnd[16]), .O(n1305) );
  ND2HHD U746 ( .I1(n1065), .I2(n1252), .O(n1068) );
  XOR2HHD U747 ( .I1(n1207), .I2(n1206), .O(n1205) );
  INVGHD U748 ( .I(n970), .O(n1207) );
  ND3CHD U749 ( .I1(n1561), .I2(n1562), .I3(n1306), .O(n1307) );
  ND2DHD U750 ( .I1(n835), .I2(n1562), .O(n836) );
  ND2DHD U751 ( .I1(n833), .I2(n1562), .O(n837) );
  XOR2HHD U752 ( .I1(n905), .I2(n906), .O(n924) );
  ND2HHD U753 ( .I1(n885), .I2(n886), .O(n905) );
  ND2HHD U754 ( .I1(n1068), .I2(n1067), .O(n1099) );
  INVCHD U755 ( .I(n1105), .O(n1007) );
  ND2DHD U756 ( .I1(n995), .I2(n994), .O(n671) );
  INVCHD U757 ( .I(n1118), .O(n1120) );
  INVCHD U758 ( .I(n1117), .O(n1121) );
  ND2DHD U759 ( .I1(n1214), .I2(n755), .O(n1254) );
  INVKHD U760 ( .I(n1137), .O(n826) );
  INVDHD U761 ( .I(n1144), .O(n1213) );
  XNR2EHD U762 ( .I1(n1252), .I2(n1253), .O(n1263) );
  ND2CHD U763 ( .I1(n1207), .I2(n1206), .O(n1208) );
  INVCHD U764 ( .I(n1233), .O(n1265) );
  ND2CHD U765 ( .I1(n1274), .I2(n1272), .O(n1278) );
  NR2CHD U766 ( .I1(n1274), .I2(n1275), .O(n711) );
  XOR2CHD U767 ( .I1(rkey_next[32]), .I2(rkey_next[13]), .O(n1453) );
  XOR2CHD U768 ( .I1(rkey_next[1]), .I2(rkey_next[36]), .O(n1411) );
  XOR2CHD U769 ( .I1(rkey_next[35]), .I2(rkey_next[0]), .O(n1497) );
  AN3CHD U770 ( .I1(n934), .I2(n1563), .I3(n933), .O(n941) );
  INVCHD U771 ( .I(rnd[23]), .O(n767) );
  ND2CHD U772 ( .I1(n937), .I2(n1305), .O(n938) );
  ND2DHD U773 ( .I1(n936), .I2(n935), .O(n939) );
  NR2BHD U774 ( .I1(rnd[5]), .I2(rnd[6]), .O(n968) );
  XOR2CHD U775 ( .I1(rnd[6]), .I2(\keyexpantion/N27 ), .O(n976) );
  ND2DHD U776 ( .I1(n801), .I2(n1568), .O(n1046) );
  AO12EHD U777 ( .B1(n974), .B2(n973), .A1(rnd[16]), .O(n993) );
  ND2HHD U778 ( .I1(n977), .I2(\keyexpantion/N27 ), .O(n995) );
  INVCKGHD U779 ( .I(n1242), .O(n882) );
  INVCHD U780 ( .I(n872), .O(n802) );
  ND2CHD U781 ( .I1(n1092), .I2(n1007), .O(n1008) );
  ND2DHD U782 ( .I1(n1005), .I2(n1105), .O(n1006) );
  ND2CHD U783 ( .I1(n1046), .I2(n1044), .O(n1075) );
  XOR2CHD U784 ( .I1(rnd[2]), .I2(rnd[7]), .O(n972) );
  ND2DHD U785 ( .I1(n1039), .I2(n1038), .O(n1074) );
  XNR2HHD U786 ( .I1(n1558), .I2(n867), .O(n898) );
  NR2EHD U787 ( .I1(n866), .I2(n878), .O(n867) );
  ND2DHD U788 ( .I1(n771), .I2(n977), .O(n952) );
  ND2DHD U789 ( .I1(n952), .I2(n984), .O(n951) );
  NR2CHD U790 ( .I1(n1027), .I2(n753), .O(n798) );
  AN2EHD U791 ( .I1(n753), .I2(n1027), .O(n758) );
  INVDHD U792 ( .I(n1112), .O(n1133) );
  ND2CHD U793 ( .I1(n1113), .I2(n1569), .O(n1116) );
  INVCHD U794 ( .I(n1000), .O(n1002) );
  OA12EHD U795 ( .B1(n983), .B2(n984), .A1(n665), .O(n1004) );
  ND2CHD U796 ( .I1(n1135), .I2(n666), .O(n665) );
  INVCHD U797 ( .I(n1032), .O(n983) );
  XNR3CHD U798 ( .I1(rnd[6]), .I2(rnd[16]), .I3(n878), .O(n870) );
  XNR2CHD U799 ( .I1(n1203), .I2(n1202), .O(n1245) );
  INVCHD U800 ( .I(n1240), .O(n1203) );
  ND2CHD U801 ( .I1(n1092), .I2(n1091), .O(n1211) );
  AN2CHD U802 ( .I1(n895), .I2(n785), .O(n618) );
  INVCHD U803 ( .I(n1245), .O(n1246) );
  INVCHD U804 ( .I(n1252), .O(n1257) );
  INVCHD U805 ( .I(n1253), .O(n1256) );
  XOR2CHD U806 ( .I1(n1251), .I2(n1250), .O(n1259) );
  OA12EHD U807 ( .B1(n1213), .B2(n1212), .A1(n1211), .O(n1249) );
  INVCHD U808 ( .I(n1210), .O(n1212) );
  OR2CHD U809 ( .I1(n1029), .I2(n1028), .O(n619) );
  ND2CHD U810 ( .I1(n1058), .I2(n1057), .O(n810) );
  INVDHD U811 ( .I(n1273), .O(n712) );
  XNR2CHD U812 ( .I1(n1265), .I2(n1264), .O(n1238) );
  INVCHD U813 ( .I(n1272), .O(n1271) );
  ND2CHD U814 ( .I1(n1579), .I2(rnd[3]), .O(n1577) );
  INVCHD U815 ( .I(n943), .O(n1316) );
  NR2BHD U816 ( .I1(rnd[26]), .I2(rnd[25]), .O(n1311) );
  NR2BHD U817 ( .I1(rnd[12]), .I2(rnd[18]), .O(n1312) );
  NR2BHD U818 ( .I1(rnd[22]), .I2(rnd[29]), .O(n1309) );
  NR2BHD U819 ( .I1(rnd[24]), .I2(rnd[23]), .O(n1310) );
  ND2CHD U820 ( .I1(n1305), .I2(n1568), .O(n1308) );
  INVDHD U821 ( .I(rnd[9]), .O(n1555) );
  AN2CHD U822 ( .I1(n1847), .I2(n1846), .O(n1848) );
  ND2CHD U823 ( .I1(n1845), .I2(key[51]), .O(n1847) );
  ND2CHD U824 ( .I1(n1807), .I2(Kin[3]), .O(n1846) );
  ND2CHD U825 ( .I1(n1852), .I2(rkey_next[3]), .O(n1853) );
  MUX2CHD U826 ( .A(n1381), .B(n1380), .S(n1379), .O(n1511) );
  ND2CHD U827 ( .I1(n1845), .I2(key[54]), .O(n1831) );
  ND2CHD U828 ( .I1(n1852), .I2(rkey_next[6]), .O(n1835) );
  ND2CHD U829 ( .I1(n1851), .I2(key[38]), .O(n1836) );
  MUX2CHD U830 ( .A(n1435), .B(n1442), .S(n1434), .O(n1823) );
  ND2CHD U831 ( .I1(n1845), .I2(key[57]), .O(n1815) );
  ND2CHD U832 ( .I1(n1852), .I2(rkey_next[9]), .O(n1819) );
  ND2CHD U833 ( .I1(n1851), .I2(key[41]), .O(n1820) );
  MUX2CHD U834 ( .A(n1424), .B(n1484), .S(n1423), .O(n1806) );
  AN2CHD U835 ( .I1(n1798), .I2(n1797), .O(n1799) );
  ND2CHD U836 ( .I1(n1845), .I2(key[60]), .O(n1798) );
  ND2CHD U837 ( .I1(n1807), .I2(Kin[12]), .O(n1797) );
  ND2CHD U838 ( .I1(n1852), .I2(rkey_next[12]), .O(n1802) );
  MUX2CHD U839 ( .A(n1391), .B(n1390), .S(n1389), .O(n1790) );
  AN2CHD U840 ( .I1(n1782), .I2(n1781), .O(n1783) );
  ND2CHD U841 ( .I1(n1845), .I2(key[63]), .O(n1782) );
  ND2CHD U842 ( .I1(n1807), .I2(Kin[15]), .O(n1781) );
  ND2CHD U843 ( .I1(n1852), .I2(rkey_next[15]), .O(n1786) );
  XNR2CHD U844 ( .I1(n1497), .I2(n1496), .O(n1774) );
  AN2CHD U845 ( .I1(n1766), .I2(n1765), .O(n1767) );
  ND2CHD U846 ( .I1(n1845), .I2(key[50]), .O(n1766) );
  ND2CHD U847 ( .I1(n1807), .I2(Kin[2]), .O(n1765) );
  ND2CHD U848 ( .I1(n1852), .I2(rkey_next[2]), .O(n1770) );
  MUX2CHD U849 ( .A(n1352), .B(n1412), .S(n1351), .O(n1758) );
  ND2CHD U850 ( .I1(n1845), .I2(key[53]), .O(n1750) );
  ND2CHD U851 ( .I1(n1852), .I2(rkey_next[5]), .O(n1754) );
  ND2CHD U852 ( .I1(n1851), .I2(key[37]), .O(n1755) );
  MUX2CHD U853 ( .A(n1444), .B(n1462), .S(n1443), .O(n1742) );
  AN2CHD U854 ( .I1(n1734), .I2(n1733), .O(n1735) );
  ND2CHD U855 ( .I1(n1845), .I2(key[56]), .O(n1734) );
  ND2CHD U856 ( .I1(n1807), .I2(Kin[8]), .O(n1733) );
  ND2CHD U857 ( .I1(n1852), .I2(rkey_next[8]), .O(n1738) );
  MUX2CHD U858 ( .A(n1487), .B(n1486), .S(n1485), .O(n1726) );
  ND2CHD U859 ( .I1(n1845), .I2(key[59]), .O(n1718) );
  ND2CHD U860 ( .I1(n1852), .I2(rkey_next[11]), .O(n1722) );
  ND2CHD U861 ( .I1(n1851), .I2(key[43]), .O(n1723) );
  MUX2CHD U862 ( .A(n1361), .B(n1400), .S(n1360), .O(n1710) );
  ND2CHD U863 ( .I1(n1845), .I2(key[62]), .O(n1702) );
  ND2CHD U864 ( .I1(n1852), .I2(rkey_next[14]), .O(n1706) );
  ND2CHD U865 ( .I1(n1851), .I2(key[46]), .O(n1707) );
  MUX2CHD U866 ( .A(n1475), .B(n1474), .S(n1473), .O(n1694) );
  ND2CHD U867 ( .I1(n1845), .I2(key[49]), .O(n1686) );
  ND2CHD U868 ( .I1(n1852), .I2(rkey_next[1]), .O(n1690) );
  ND2CHD U869 ( .I1(n1851), .I2(key[33]), .O(n1691) );
  XNR2CHD U870 ( .I1(n1414), .I2(n1413), .O(n1682) );
  MUX2CHD U871 ( .A(rkey[1]), .B(n1689), .S(n1412), .O(n1413) );
  ND2CHD U872 ( .I1(n1845), .I2(key[52]), .O(n1674) );
  ND2CHD U873 ( .I1(n1852), .I2(rkey_next[4]), .O(n1678) );
  ND2CHD U874 ( .I1(n1851), .I2(key[36]), .O(n1679) );
  MUX2CHD U875 ( .A(n1465), .B(n1464), .S(n1463), .O(n1506) );
  AN2CHD U876 ( .I1(n1661), .I2(n1660), .O(n1662) );
  ND2CHD U877 ( .I1(n1845), .I2(key[55]), .O(n1661) );
  ND2CHD U878 ( .I1(n1807), .I2(Kin[7]), .O(n1660) );
  ND2CHD U879 ( .I1(n1852), .I2(rkey_next[7]), .O(n1665) );
  MUX2CHD U880 ( .A(n1371), .B(n1433), .S(n1370), .O(n1653) );
  ND2CHD U881 ( .I1(n1845), .I2(key[58]), .O(n1645) );
  ND2CHD U882 ( .I1(n1852), .I2(rkey_next[10]), .O(n1649) );
  ND2CHD U883 ( .I1(n1851), .I2(key[42]), .O(n1650) );
  MUX2CHD U884 ( .A(n1402), .B(n1422), .S(n1401), .O(n1637) );
  AN2CHD U885 ( .I1(n1629), .I2(n1628), .O(n1630) );
  ND2CHD U886 ( .I1(n1845), .I2(key[61]), .O(n1629) );
  ND2CHD U887 ( .I1(n1807), .I2(Kin[13]), .O(n1628) );
  ND2CHD U888 ( .I1(n1852), .I2(rkey_next[13]), .O(n1633) );
  ND2CHD U889 ( .I1(n1807), .I2(Kin[29]), .O(n1624) );
  XNR2CHD U890 ( .I1(n1453), .I2(n1452), .O(n1621) );
  MUX2CHD U891 ( .A(rkey[13]), .B(n1632), .S(n1474), .O(n1452) );
  XNR3CHD U892 ( .I1(rkey[0]), .I2(n1411), .I3(n1497), .O(n1548) );
  ND2CHD U893 ( .I1(n1807), .I2(Kin[48]), .O(n1587) );
  INVCHD U894 ( .I(n1852), .O(n1551) );
  INVCHD U895 ( .I(n915), .O(n854) );
  ND2CHD U896 ( .I1(n844), .I2(n843), .O(n846) );
  INVCHD U897 ( .I(rnd[4]), .O(n843) );
  INVDHD U898 ( .I(n990), .O(n740) );
  ND2DHD U899 ( .I1(n990), .I2(n788), .O(n739) );
  NR2EHD U900 ( .I1(n869), .I2(n868), .O(n973) );
  INVCHD U901 ( .I(n1039), .O(n887) );
  INVDHD U902 ( .I(n1251), .O(n889) );
  ND2CHD U903 ( .I1(n969), .I2(n1579), .O(n1037) );
  ND2CHD U904 ( .I1(n1013), .I2(n863), .O(n874) );
  NR2BHD U905 ( .I1(n828), .I2(n830), .O(n829) );
  ND2CHD U906 ( .I1(n943), .I2(rnd[20]), .O(n828) );
  INVCHD U907 ( .I(n830), .O(n831) );
  NR2BHD U908 ( .I1(rnd[8]), .I2(rnd[7]), .O(n853) );
  AN2CHD U909 ( .I1(n941), .I2(n767), .O(n625) );
  ND2CHD U910 ( .I1(n745), .I2(n1579), .O(n1105) );
  INVCHD U911 ( .I(n985), .O(n986) );
  INVCHD U912 ( .I(n1044), .O(n1090) );
  XNR2CHD U913 ( .I1(n1579), .I2(n981), .O(n1108) );
  XOR2CHD U914 ( .I1(rnd[13]), .I2(rnd[3]), .O(n981) );
  ND2DHD U915 ( .I1(n823), .I2(n790), .O(n789) );
  AN2CHD U916 ( .I1(n934), .I2(n1562), .O(n790) );
  INVCHD U917 ( .I(n822), .O(n823) );
  ND2DHD U918 ( .I1(n786), .I2(n974), .O(n751) );
  AN2CHD U919 ( .I1(n974), .I2(n824), .O(n749) );
  INVCHD U920 ( .I(n1073), .O(n1098) );
  ND2CHD U921 ( .I1(n1071), .I2(n1070), .O(n1100) );
  ND2CHD U922 ( .I1(n1069), .I2(rnd[14]), .O(n1070) );
  INVCHD U923 ( .I(n993), .O(n992) );
  AN2CHD U924 ( .I1(n1106), .I2(n1105), .O(n1112) );
  ND2DHD U925 ( .I1(n1136), .I2(rnd[12]), .O(n1106) );
  AN2CHD U926 ( .I1(n1001), .I2(n998), .O(n622) );
  ND2DHD U927 ( .I1(n1052), .I2(n1054), .O(n697) );
  INVCHD U928 ( .I(n1076), .O(n1049) );
  ND2CHD U929 ( .I1(n1077), .I2(n1075), .O(n1050) );
  ND2DHD U930 ( .I1(n673), .I2(n669), .O(n698) );
  ND2CHD U931 ( .I1(n884), .I2(rnd[30]), .O(n885) );
  ND2CHD U932 ( .I1(n1039), .I2(n1045), .O(n891) );
  ND2CHD U933 ( .I1(n887), .I2(n1090), .O(n888) );
  ND2DHD U934 ( .I1(n1140), .I2(n912), .O(n911) );
  XNR2CHD U935 ( .I1(rnd[5]), .I2(n1037), .O(n1038) );
  NR2BHD U936 ( .I1(rnd[14]), .I2(n869), .O(n839) );
  ND2CHD U937 ( .I1(n853), .I2(n914), .O(n879) );
  INVCHD U938 ( .I(n910), .O(n851) );
  XNR2HHD U939 ( .I1(rnd[8]), .I2(n944), .O(n982) );
  NR2CHD U940 ( .I1(n1014), .I2(n1033), .O(n1015) );
  XOR2EHD U941 ( .I1(rnd[28]), .I2(n949), .O(n970) );
  ND2DHD U942 ( .I1(n768), .I2(n948), .O(n949) );
  NR2CHD U943 ( .I1(n947), .I2(n1033), .O(n948) );
  XNR2CHD U944 ( .I1(rnd[7]), .I2(n971), .O(n950) );
  ND2DHD U945 ( .I1(n691), .I2(n1023), .O(n690) );
  XNR2CHD U946 ( .I1(rnd[31]), .I2(n1061), .O(n1064) );
  ND2DHD U947 ( .I1(n702), .I2(n1100), .O(n701) );
  ND3CHD U948 ( .I1(n1068), .I2(n1067), .I3(n703), .O(n702) );
  INVCKGHD U949 ( .I(n1111), .O(n1131) );
  OR2CHD U950 ( .I1(n754), .I2(n982), .O(n621) );
  INVCHD U951 ( .I(n1107), .O(n754) );
  NR2CHD U952 ( .I1(n788), .I2(n789), .O(n787) );
  ND2DHD U953 ( .I1(n1073), .I2(rnd[25]), .O(n719) );
  INVDHD U954 ( .I(n1078), .O(n645) );
  INVDHD U955 ( .I(n1024), .O(n893) );
  ND2CHD U956 ( .I1(n903), .I2(n902), .O(n904) );
  INVCHD U957 ( .I(n906), .O(n903) );
  INVCHD U958 ( .I(n905), .O(n902) );
  XNR3CHD U959 ( .I1(n1061), .I2(n897), .I3(n896), .O(n923) );
  ND2CHD U960 ( .I1(n906), .I2(n905), .O(n925) );
  ND2DHD U961 ( .I1(n913), .I2(n991), .O(n638) );
  ND2DHD U962 ( .I1(n911), .I2(n989), .O(n637) );
  INVCHD U963 ( .I(n912), .O(n913) );
  ND3CHD U964 ( .I1(n974), .I2(n824), .I3(n1350), .O(n678) );
  XNR2CHD U965 ( .I1(n982), .I2(n1214), .O(n1210) );
  MAO222CHD U966 ( .A1(n1135), .B1(n950), .C1(rnd[17]), .O(n1206) );
  ND2CHD U967 ( .I1(n1110), .I2(n953), .O(n954) );
  INVCHD U968 ( .I(n952), .O(n953) );
  XOR2EHD U969 ( .I1(n1205), .I2(n1204), .O(n1199) );
  INVDHD U970 ( .I(n1159), .O(n687) );
  ND2DHD U971 ( .I1(n1165), .I2(n733), .O(n686) );
  ND2CHD U972 ( .I1(n1163), .I2(n1162), .O(n1165) );
  INVCHD U973 ( .I(n1161), .O(n1162) );
  XNR2EHD U974 ( .I1(n923), .I2(n924), .O(n1167) );
  ND2DHD U975 ( .I1(n1166), .I2(\keyexpantion/N27 ), .O(n1171) );
  ND2DHD U976 ( .I1(n806), .I2(n805), .O(n1166) );
  ND2CHD U977 ( .I1(n1102), .I2(n1101), .O(n1103) );
  ND2CHD U978 ( .I1(n1127), .I2(n1128), .O(n1104) );
  XOR2CHD U979 ( .I1(n1134), .I2(n616), .O(n1147) );
  MAO222CHD U980 ( .A1(n1131), .B1(n1130), .C1(n1110), .O(n1134) );
  XOR2CHD U981 ( .I1(n1133), .I2(n1132), .O(n616) );
  XOR2CHD U982 ( .I1(n1213), .I2(rnd[28]), .O(n1145) );
  MAO222CHD U983 ( .A1(n1143), .B1(n1142), .C1(n1141), .O(n1146) );
  XNR2CHD U984 ( .I1(n1136), .I2(n1135), .O(n1142) );
  MAO222CHD U985 ( .A1(n1140), .B1(n1139), .C1(n1138), .O(n1141) );
  ND2CHD U986 ( .I1(n1137), .I2(\keyexpantion/N26 ), .O(n1139) );
  OA12EHD U987 ( .B1(n1126), .B2(n1129), .A1(n1125), .O(n1149) );
  INVCHD U988 ( .I(n1122), .O(n1124) );
  OR2CHD U989 ( .I1(n1004), .I2(n1003), .O(n815) );
  ND2CHD U990 ( .I1(n900), .I2(n899), .O(n901) );
  INVCHD U991 ( .I(n956), .O(n929) );
  ND2DHD U992 ( .I1(n926), .I2(n925), .O(n962) );
  ND2CHD U993 ( .I1(n924), .I2(n923), .O(n926) );
  OA12EHD U994 ( .B1(n929), .B2(n961), .A1(n960), .O(n1195) );
  ND2CHD U995 ( .I1(n959), .I2(n958), .O(n960) );
  INVCHD U996 ( .I(n957), .O(n958) );
  XNR2CHD U997 ( .I1(rnd[3]), .I2(rnd[2]), .O(n1190) );
  INVCHD U998 ( .I(n716), .O(n715) );
  XNR3CHD U999 ( .I1(n1262), .I2(n1261), .I3(n1260), .O(n1267) );
  XOR2CHD U1000 ( .I1(n1244), .I2(n1243), .O(n1262) );
  XNR2CHD U1001 ( .I1(n1234), .I2(n1233), .O(n1217) );
  INVCHD U1002 ( .I(n1235), .O(n1237) );
  ND2HHD U1003 ( .I1(n775), .I2(n774), .O(n1177) );
  INVDHD U1004 ( .I(n1169), .O(n774) );
  INVDHD U1005 ( .I(n1168), .O(n775) );
  INVCHD U1006 ( .I(n1183), .O(n1175) );
  INVDHD U1007 ( .I(n964), .O(n967) );
  NR2BHD U1008 ( .I1(n657), .I2(n1059), .O(n811) );
  ND2HHD U1009 ( .I1(n965), .I2(n964), .O(n1230) );
  INVCHD U1010 ( .I(n1285), .O(n1280) );
  INVCHD U1011 ( .I(sel), .O(n1294) );
  ND3CHD U1012 ( .I1(n712), .I2(n1277), .I3(n711), .O(n710) );
  INVCHD U1013 ( .I(Krdy), .O(n1327) );
  XOR2CHD U1014 ( .I1(n818), .I2(n1548), .O(n626) );
  OR2CHD U1015 ( .I1(Drdy), .I2(n1297), .O(n1298) );
  INVCHD U1016 ( .I(rnd[30]), .O(n1568) );
  INVCHD U1017 ( .I(rnd[29]), .O(n1569) );
  INVCHD U1018 ( .I(rnd[26]), .O(n1565) );
  INVDHD U1019 ( .I(rnd[25]), .O(n1566) );
  INVDHD U1020 ( .I(rnd[24]), .O(n1564) );
  INVDHD U1021 ( .I(rnd[22]), .O(n1563) );
  INVCHD U1022 ( .I(rnd[21]), .O(n788) );
  INVDHD U1023 ( .I(rnd[18]), .O(n1560) );
  INVDHD U1024 ( .I(rnd[16]), .O(n909) );
  INVCHD U1025 ( .I(rnd[12]), .O(n1557) );
  INVDHD U1026 ( .I(rnd[11]), .O(n1558) );
  INVDHD U1027 ( .I(rnd[10]), .O(n1556) );
  INVCHD U1028 ( .I(Drdy), .O(n1348) );
  ND2CHD U1029 ( .I1(n1807), .I2(Kin[35]), .O(n1613) );
  ND2CHD U1030 ( .I1(n1807), .I2(Kin[38]), .O(n1607) );
  ND2CHD U1031 ( .I1(n1807), .I2(Kin[41]), .O(n1601) );
  ND2CHD U1032 ( .I1(n1807), .I2(Kin[44]), .O(n1595) );
  ND2CHD U1033 ( .I1(n1807), .I2(Kin[47]), .O(n1589) );
  ND2CHD U1034 ( .I1(n1807), .I2(Kin[34]), .O(n1615) );
  ND2CHD U1035 ( .I1(n1807), .I2(Kin[37]), .O(n1609) );
  ND2CHD U1036 ( .I1(n1807), .I2(Kin[40]), .O(n1603) );
  ND2CHD U1037 ( .I1(n1807), .I2(Kin[43]), .O(n1597) );
  ND2CHD U1038 ( .I1(n1807), .I2(Kin[46]), .O(n1591) );
  ND2CHD U1039 ( .I1(n1807), .I2(Kin[33]), .O(n1617) );
  ND2CHD U1040 ( .I1(n1807), .I2(Kin[36]), .O(n1611) );
  ND2CHD U1041 ( .I1(n1807), .I2(Kin[39]), .O(n1605) );
  ND2CHD U1042 ( .I1(n1807), .I2(Kin[42]), .O(n1599) );
  ND2CHD U1043 ( .I1(n1807), .I2(Kin[45]), .O(n1593) );
  NR2BHD U1044 ( .I1(n1578), .I2(n1329), .O(n1330) );
  ND2CHD U1045 ( .I1(n1807), .I2(Kin[32]), .O(n1619) );
  NR2BHD U1046 ( .I1(Drdy), .I2(rnd[13]), .O(n1301) );
  NR2BHD U1047 ( .I1(rnd[21]), .I2(rnd[27]), .O(n1304) );
  NR2BHD U1048 ( .I1(n1316), .I2(n1315), .O(n1317) );
  ND2CHD U1049 ( .I1(n1326), .I2(n1325), .O(n611) );
  AO222CHD U1050 ( .A1(n1571), .A2(Dout[6]), .B1(n1573), .B2(Din[6]), .C1(
        n1572), .C2(dat_next[6]), .O(n510) );
  ND2CHD U1051 ( .I1(n1441), .I2(n1440), .O(n494) );
  AO222CHD U1052 ( .A1(n1571), .A2(Dout[5]), .B1(n1573), .B2(Din[5]), .C1(
        n1572), .C2(dat_next[5]), .O(n511) );
  ND2CHD U1053 ( .I1(n1451), .I2(n1450), .O(n495) );
  AO222CHD U1054 ( .A1(n1571), .A2(Dout[13]), .B1(n1573), .B2(Din[13]), .C1(
        n1572), .C2(dat_next[13]), .O(n503) );
  ND2CHD U1055 ( .I1(n1461), .I2(n1460), .O(n487) );
  AO222CHD U1056 ( .A1(n1571), .A2(Dout[4]), .B1(n1573), .B2(Din[4]), .C1(
        n1572), .C2(dat_next[4]), .O(n512) );
  ND2CHD U1057 ( .I1(n1472), .I2(n1471), .O(n496) );
  AO222CHD U1058 ( .A1(n1571), .A2(Dout[3]), .B1(n1573), .B2(Din[3]), .C1(
        n1572), .C2(dat_next[3]), .O(n513) );
  ND2CHD U1059 ( .I1(n1388), .I2(n1387), .O(n497) );
  AO222CHD U1060 ( .A1(n1571), .A2(Dout[11]), .B1(n1573), .B2(Din[11]), .C1(
        n1572), .C2(dat_next[11]), .O(n505) );
  ND2CHD U1061 ( .I1(n1369), .I2(n1368), .O(n489) );
  AO222CHD U1062 ( .A1(n1571), .A2(Dout[2]), .B1(n1573), .B2(Din[2]), .C1(
        n1572), .C2(dat_next[2]), .O(n514) );
  ND2CHD U1063 ( .I1(n1359), .I2(n1358), .O(n498) );
  AO222CHD U1064 ( .A1(n1571), .A2(Dout[1]), .B1(n1573), .B2(Din[1]), .C1(
        n1572), .C2(dat_next[1]), .O(n515) );
  ND2CHD U1065 ( .I1(n1421), .I2(n1420), .O(n499) );
  AO222CHD U1066 ( .A1(n1571), .A2(Dout[9]), .B1(n1573), .B2(Din[9]), .C1(
        n1572), .C2(dat_next[9]), .O(n507) );
  ND2CHD U1067 ( .I1(n1432), .I2(n1431), .O(n491) );
  AO222CHD U1068 ( .A1(n1571), .A2(Dout[7]), .B1(n1573), .B2(Din[7]), .C1(
        n1572), .C2(dat_next[7]), .O(n509) );
  ND2CHD U1069 ( .I1(n1378), .I2(n1377), .O(n493) );
  AO222CHD U1070 ( .A1(n1571), .A2(Dout[15]), .B1(n1573), .B2(Din[15]), .C1(
        n1572), .C2(dat_next[15]), .O(n501) );
  ND2CHD U1071 ( .I1(n1505), .I2(n1504), .O(n484) );
  AO222CHD U1072 ( .A1(n1571), .A2(Dout[14]), .B1(n1573), .B2(Din[14]), .C1(
        n1572), .C2(dat_next[14]), .O(n502) );
  ND2CHD U1073 ( .I1(n1483), .I2(n1482), .O(n486) );
  AO222CHD U1074 ( .A1(n1571), .A2(Dout[12]), .B1(n1573), .B2(Din[12]), .C1(
        n1572), .C2(dat_next[12]), .O(n504) );
  ND2CHD U1075 ( .I1(n1399), .I2(n1398), .O(n488) );
  AO222CHD U1076 ( .A1(n1571), .A2(Dout[10]), .B1(n1573), .B2(Din[10]), .C1(
        n1572), .C2(dat_next[10]), .O(n506) );
  ND2CHD U1077 ( .I1(n1410), .I2(n1409), .O(n490) );
  AO222CHD U1078 ( .A1(n1571), .A2(Dout[8]), .B1(n1573), .B2(Din[8]), .C1(
        n1572), .C2(dat_next[8]), .O(n508) );
  ND2CHD U1079 ( .I1(n1494), .I2(n1493), .O(n492) );
  ND2CHD U1080 ( .I1(n1572), .I2(dat_next[0]), .O(n1575) );
  ND2CHD U1081 ( .I1(n1571), .I2(Dout[0]), .O(n1576) );
  MUX2CHD U1082 ( .A(key[0]), .B(Kin[0]), .S(n1807), .O(n517) );
  MUX2CHD U1083 ( .A(key[1]), .B(Kin[1]), .S(n1807), .O(n518) );
  MUX2CHD U1084 ( .A(key[2]), .B(Kin[2]), .S(n1807), .O(n519) );
  MUX2CHD U1085 ( .A(key[3]), .B(Kin[3]), .S(n1807), .O(n520) );
  MUX2CHD U1086 ( .A(key[4]), .B(Kin[4]), .S(n1807), .O(n521) );
  MUX2CHD U1087 ( .A(key[5]), .B(Kin[5]), .S(n1807), .O(n522) );
  MUX2CHD U1088 ( .A(key[6]), .B(Kin[6]), .S(n1807), .O(n523) );
  MUX2CHD U1089 ( .A(key[7]), .B(Kin[7]), .S(n1807), .O(n524) );
  MUX2CHD U1090 ( .A(key[8]), .B(Kin[8]), .S(n1807), .O(n525) );
  MUX2CHD U1091 ( .A(key[9]), .B(Kin[9]), .S(n1807), .O(n526) );
  MUX2CHD U1092 ( .A(key[10]), .B(Kin[10]), .S(n1807), .O(n527) );
  MUX2CHD U1093 ( .A(key[11]), .B(Kin[11]), .S(n1807), .O(n528) );
  MUX2CHD U1094 ( .A(key[12]), .B(Kin[12]), .S(n1807), .O(n529) );
  MUX2CHD U1095 ( .A(key[13]), .B(Kin[13]), .S(n1807), .O(n530) );
  MUX2CHD U1096 ( .A(key[14]), .B(Kin[14]), .S(n1807), .O(n531) );
  MUX2CHD U1097 ( .A(key[15]), .B(Kin[15]), .S(n1807), .O(n532) );
  MUX2CHD U1098 ( .A(key[16]), .B(Kin[16]), .S(n1807), .O(n533) );
  MUX2CHD U1099 ( .A(key[17]), .B(Kin[17]), .S(n1807), .O(n534) );
  MUX2CHD U1100 ( .A(key[18]), .B(Kin[18]), .S(n1807), .O(n535) );
  MUX2CHD U1101 ( .A(key[19]), .B(Kin[19]), .S(n1807), .O(n536) );
  MUX2CHD U1102 ( .A(key[20]), .B(Kin[20]), .S(n1807), .O(n537) );
  MUX2CHD U1103 ( .A(key[21]), .B(Kin[21]), .S(n1807), .O(n538) );
  MUX2CHD U1104 ( .A(key[22]), .B(Kin[22]), .S(n1807), .O(n539) );
  MUX2CHD U1105 ( .A(key[23]), .B(Kin[23]), .S(n1807), .O(n540) );
  MUX2CHD U1106 ( .A(key[24]), .B(Kin[24]), .S(n1807), .O(n541) );
  MUX2CHD U1107 ( .A(key[25]), .B(Kin[25]), .S(n1807), .O(n542) );
  MUX2CHD U1108 ( .A(key[26]), .B(Kin[26]), .S(n1807), .O(n543) );
  MUX2CHD U1109 ( .A(key[27]), .B(Kin[27]), .S(n1807), .O(n544) );
  MUX2CHD U1110 ( .A(key[28]), .B(Kin[28]), .S(n1807), .O(n545) );
  MUX2CHD U1111 ( .A(key[29]), .B(Kin[29]), .S(n1807), .O(n546) );
  MUX2CHD U1112 ( .A(key[30]), .B(Kin[30]), .S(n1807), .O(n547) );
  MUX2CHD U1113 ( .A(key[31]), .B(Kin[31]), .S(n1807), .O(n548) );
  MUX2CHD U1114 ( .A(key[49]), .B(Kin[49]), .S(n1807), .O(n566) );
  MUX2CHD U1115 ( .A(key[50]), .B(Kin[50]), .S(n1807), .O(n567) );
  MUX2CHD U1116 ( .A(key[51]), .B(Kin[51]), .S(n1807), .O(n568) );
  MUX2CHD U1117 ( .A(key[52]), .B(Kin[52]), .S(n1807), .O(n569) );
  MUX2CHD U1118 ( .A(key[53]), .B(Kin[53]), .S(n1807), .O(n570) );
  MUX2CHD U1119 ( .A(key[54]), .B(Kin[54]), .S(n1807), .O(n571) );
  MUX2CHD U1120 ( .A(key[55]), .B(Kin[55]), .S(n1807), .O(n572) );
  MUX2CHD U1121 ( .A(key[56]), .B(Kin[56]), .S(n1807), .O(n573) );
  MUX2CHD U1122 ( .A(key[57]), .B(Kin[57]), .S(n1807), .O(n574) );
  MUX2CHD U1123 ( .A(key[58]), .B(Kin[58]), .S(n1807), .O(n575) );
  MUX2CHD U1124 ( .A(key[59]), .B(Kin[59]), .S(n1807), .O(n576) );
  MUX2CHD U1125 ( .A(key[60]), .B(Kin[60]), .S(n1807), .O(n577) );
  MUX2CHD U1126 ( .A(key[61]), .B(Kin[61]), .S(n1807), .O(n578) );
  MUX2CHD U1127 ( .A(key[62]), .B(Kin[62]), .S(n1807), .O(n579) );
  MUX2CHD U1128 ( .A(key[63]), .B(Kin[63]), .S(n1807), .O(n580) );
  MUX2CHD U1129 ( .A(rnd[30]), .B(rnd[31]), .S(n1570), .O(n612) );
  MUX2CHD U1130 ( .A(rnd[27]), .B(rnd[28]), .S(n1570), .O(n583) );
  MUX2CHD U1131 ( .A(rnd[26]), .B(rnd[27]), .S(n1570), .O(n584) );
  MUX2CHD U1132 ( .A(rnd[23]), .B(rnd[24]), .S(n1570), .O(n587) );
  MUX2CHD U1133 ( .A(rnd[22]), .B(rnd[23]), .S(n1570), .O(n588) );
  MXL2CHD U1134 ( .A(n1562), .B(n788), .S(n1570), .OB(n590) );
  MUX2CHD U1135 ( .A(rnd[17]), .B(rnd[18]), .S(n1570), .O(n593) );
  MUX2CHD U1136 ( .A(rnd[16]), .B(rnd[17]), .S(n1570), .O(n594) );
  MUX2CHD U1137 ( .A(rnd[13]), .B(rnd[14]), .S(n1570), .O(n597) );
  MUX2CHD U1138 ( .A(rnd[12]), .B(rnd[13]), .S(n1570), .O(n598) );
  INVCHD U1139 ( .I(rnd[8]), .O(n1554) );
  MUX2CHD U1140 ( .A(rnd[7]), .B(rnd[8]), .S(n1570), .O(n603) );
  MUX2CHD U1141 ( .A(rnd[6]), .B(rnd[7]), .S(n1570), .O(n604) );
  MUX2CHD U1142 ( .A(rnd[5]), .B(rnd[6]), .S(n1570), .O(n605) );
  MUX2CHD U1143 ( .A(rnd[4]), .B(rnd[5]), .S(n1570), .O(n606) );
  MUX2CHD U1144 ( .A(rnd[3]), .B(rnd[4]), .S(n1570), .O(n607) );
  MUX2CHD U1145 ( .A(rnd[2]), .B(rnd[3]), .S(n1570), .O(n608) );
  AN2CHD U1146 ( .I1(n1854), .I2(n1853), .O(n1855) );
  ND2CHD U1147 ( .I1(n1851), .I2(key[35]), .O(n1854) );
  AN2CHD U1148 ( .I1(n1840), .I2(n1839), .O(n1841) );
  ND2CHD U1149 ( .I1(n1852), .I2(rkey_next[19]), .O(n1840) );
  ND2CHD U1150 ( .I1(n1807), .I2(Kin[19]), .O(n1839) );
  ND2CHD U1151 ( .I1(n1335), .I2(n1613), .O(n418) );
  AN2CHD U1152 ( .I1(n1334), .I2(n1333), .O(n1335) );
  ND2CHD U1153 ( .I1(rkey_next[19]), .I2(n1584), .O(n1333) );
  ND2CHD U1154 ( .I1(n1852), .I2(rkey_next[35]), .O(n1334) );
  ND2CHD U1155 ( .I1(n1513), .I2(n1512), .O(n419) );
  ND2CHD U1156 ( .I1(n1511), .I2(n1852), .O(n1513) );
  AN2CHD U1157 ( .I1(n1836), .I2(n1835), .O(n1837) );
  AN2CHD U1158 ( .I1(n1831), .I2(n1830), .O(n1832) );
  AN2CHD U1159 ( .I1(n1827), .I2(n1826), .O(n1828) );
  ND2CHD U1160 ( .I1(n1807), .I2(Kin[22]), .O(n1826) );
  ND2CHD U1161 ( .I1(n1852), .I2(rkey_next[22]), .O(n1827) );
  ND2CHD U1162 ( .I1(n1528), .I2(n1607), .O(n422) );
  AN2CHD U1163 ( .I1(n1527), .I2(n1526), .O(n1528) );
  ND2CHD U1164 ( .I1(rkey_next[22]), .I2(n1584), .O(n1526) );
  ND2CHD U1165 ( .I1(n1852), .I2(rkey_next[38]), .O(n1527) );
  AN2CHD U1166 ( .I1(n1820), .I2(n1819), .O(n1821) );
  AN2CHD U1167 ( .I1(n1815), .I2(n1814), .O(n1816) );
  AN2CHD U1168 ( .I1(n1811), .I2(n1810), .O(n1812) );
  ND2CHD U1169 ( .I1(n1852), .I2(rkey_next[25]), .O(n1811) );
  ND2CHD U1170 ( .I1(n1807), .I2(Kin[25]), .O(n1810) );
  ND2CHD U1171 ( .I1(n1534), .I2(n1601), .O(n426) );
  AN2CHD U1172 ( .I1(n1533), .I2(n1532), .O(n1534) );
  ND2CHD U1173 ( .I1(rkey_next[25]), .I2(n1584), .O(n1532) );
  ND2CHD U1174 ( .I1(n1852), .I2(rkey_next[41]), .O(n1533) );
  AN2CHD U1175 ( .I1(n1803), .I2(n1802), .O(n1804) );
  ND2CHD U1176 ( .I1(n1851), .I2(key[44]), .O(n1803) );
  AN2CHD U1177 ( .I1(n1794), .I2(n1793), .O(n1795) );
  ND2CHD U1178 ( .I1(n1807), .I2(Kin[28]), .O(n1793) );
  ND2CHD U1179 ( .I1(n1852), .I2(rkey_next[28]), .O(n1794) );
  ND2CHD U1180 ( .I1(n1341), .I2(n1595), .O(n430) );
  AN2CHD U1181 ( .I1(n1340), .I2(n1339), .O(n1341) );
  ND2CHD U1182 ( .I1(rkey_next[28]), .I2(n1584), .O(n1339) );
  ND2CHD U1183 ( .I1(n1852), .I2(rkey_next[44]), .O(n1340) );
  AN2CHD U1184 ( .I1(n1787), .I2(n1786), .O(n1788) );
  ND2CHD U1185 ( .I1(n1851), .I2(key[47]), .O(n1787) );
  AN2CHD U1186 ( .I1(n1778), .I2(n1777), .O(n1779) );
  ND2CHD U1187 ( .I1(n1807), .I2(Kin[31]), .O(n1777) );
  ND2CHD U1188 ( .I1(n1852), .I2(rkey_next[31]), .O(n1778) );
  ND2CHD U1189 ( .I1(n1531), .I2(n1589), .O(n434) );
  AN2CHD U1190 ( .I1(n1530), .I2(n1529), .O(n1531) );
  ND2CHD U1191 ( .I1(rkey_next[31]), .I2(n1584), .O(n1529) );
  ND2CHD U1192 ( .I1(n1852), .I2(rkey_next[47]), .O(n1530) );
  AN2CHD U1193 ( .I1(n1771), .I2(n1770), .O(n1772) );
  ND2CHD U1194 ( .I1(n1851), .I2(key[34]), .O(n1771) );
  AN2CHD U1195 ( .I1(n1762), .I2(n1761), .O(n1763) );
  ND2CHD U1196 ( .I1(n1807), .I2(Kin[18]), .O(n1761) );
  ND2CHD U1197 ( .I1(n1852), .I2(rkey_next[18]), .O(n1762) );
  ND2CHD U1198 ( .I1(n1338), .I2(n1615), .O(n438) );
  AN2CHD U1199 ( .I1(n1337), .I2(n1336), .O(n1338) );
  ND2CHD U1200 ( .I1(rkey_next[18]), .I2(n1584), .O(n1336) );
  ND2CHD U1201 ( .I1(n1852), .I2(rkey_next[34]), .O(n1337) );
  AN2CHD U1202 ( .I1(n1755), .I2(n1754), .O(n1756) );
  AN2CHD U1203 ( .I1(n1750), .I2(n1749), .O(n1751) );
  AN2CHD U1204 ( .I1(n1746), .I2(n1745), .O(n1747) );
  ND2CHD U1205 ( .I1(n1807), .I2(Kin[21]), .O(n1745) );
  ND2CHD U1206 ( .I1(n1852), .I2(rkey_next[21]), .O(n1746) );
  ND2CHD U1207 ( .I1(n1522), .I2(n1609), .O(n442) );
  AN2CHD U1208 ( .I1(n1521), .I2(n1520), .O(n1522) );
  ND2CHD U1209 ( .I1(rkey_next[21]), .I2(n1584), .O(n1520) );
  ND2CHD U1210 ( .I1(n1852), .I2(rkey_next[37]), .O(n1521) );
  AN2CHD U1211 ( .I1(n1739), .I2(n1738), .O(n1740) );
  ND2CHD U1212 ( .I1(n1851), .I2(key[40]), .O(n1739) );
  AN2CHD U1213 ( .I1(n1730), .I2(n1729), .O(n1731) );
  ND2CHD U1214 ( .I1(n1852), .I2(rkey_next[24]), .O(n1730) );
  ND2CHD U1215 ( .I1(n1807), .I2(Kin[24]), .O(n1729) );
  ND2CHD U1216 ( .I1(n1537), .I2(n1603), .O(n446) );
  AN2CHD U1217 ( .I1(n1536), .I2(n1535), .O(n1537) );
  ND2CHD U1218 ( .I1(rkey_next[24]), .I2(n1584), .O(n1535) );
  ND2CHD U1219 ( .I1(n1852), .I2(rkey_next[40]), .O(n1536) );
  AN2CHD U1220 ( .I1(n1723), .I2(n1722), .O(n1724) );
  AN2CHD U1221 ( .I1(n1718), .I2(n1717), .O(n1719) );
  AN2CHD U1222 ( .I1(n1714), .I2(n1713), .O(n1715) );
  ND2CHD U1223 ( .I1(n1807), .I2(Kin[27]), .O(n1713) );
  ND2CHD U1224 ( .I1(n1852), .I2(rkey_next[27]), .O(n1714) );
  ND2CHD U1225 ( .I1(n1344), .I2(n1597), .O(n450) );
  AN2CHD U1226 ( .I1(n1343), .I2(n1342), .O(n1344) );
  ND2CHD U1227 ( .I1(rkey_next[27]), .I2(n1584), .O(n1342) );
  ND2CHD U1228 ( .I1(n1852), .I2(rkey_next[43]), .O(n1343) );
  AN2CHD U1229 ( .I1(n1707), .I2(n1706), .O(n1708) );
  AN2CHD U1230 ( .I1(n1702), .I2(n1701), .O(n1703) );
  AN2CHD U1231 ( .I1(n1698), .I2(n1697), .O(n1699) );
  ND2CHD U1232 ( .I1(n1852), .I2(rkey_next[30]), .O(n1698) );
  ND2CHD U1233 ( .I1(n1807), .I2(Kin[30]), .O(n1697) );
  ND2CHD U1234 ( .I1(n1519), .I2(n1591), .O(n454) );
  AN2CHD U1235 ( .I1(n1518), .I2(n1517), .O(n1519) );
  ND2CHD U1236 ( .I1(rkey_next[30]), .I2(n1584), .O(n1517) );
  ND2CHD U1237 ( .I1(n1852), .I2(rkey_next[46]), .O(n1518) );
  AN2CHD U1238 ( .I1(n1691), .I2(n1690), .O(n1692) );
  AN2CHD U1239 ( .I1(n1686), .I2(n1685), .O(n1687) );
  ND2CHD U1240 ( .I1(n1332), .I2(n1331), .O(n457) );
  ND2CHD U1241 ( .I1(n1852), .I2(rkey_next[17]), .O(n1332) );
  ND2CHD U1242 ( .I1(n1525), .I2(n1617), .O(n458) );
  AN2CHD U1243 ( .I1(n1524), .I2(n1523), .O(n1525) );
  ND2CHD U1244 ( .I1(rkey_next[17]), .I2(n1584), .O(n1523) );
  ND2CHD U1245 ( .I1(n1852), .I2(rkey_next[33]), .O(n1524) );
  AN2CHD U1246 ( .I1(n1679), .I2(n1678), .O(n1680) );
  AN2CHD U1247 ( .I1(n1674), .I2(n1673), .O(n1675) );
  AN2CHD U1248 ( .I1(n1670), .I2(n1669), .O(n1671) );
  ND2CHD U1249 ( .I1(n1852), .I2(rkey_next[20]), .O(n1670) );
  ND2CHD U1250 ( .I1(n1807), .I2(Kin[20]), .O(n1669) );
  ND2CHD U1251 ( .I1(n1543), .I2(n1611), .O(n462) );
  AN2CHD U1252 ( .I1(n1542), .I2(n1541), .O(n1543) );
  ND2CHD U1253 ( .I1(rkey_next[20]), .I2(n1584), .O(n1541) );
  ND2CHD U1254 ( .I1(n1852), .I2(rkey_next[36]), .O(n1542) );
  ND2CHD U1255 ( .I1(n1508), .I2(n1507), .O(n463) );
  ND2CHD U1256 ( .I1(n1506), .I2(n1852), .O(n1508) );
  AN2CHD U1257 ( .I1(n1666), .I2(n1665), .O(n1667) );
  ND2CHD U1258 ( .I1(n1851), .I2(key[39]), .O(n1666) );
  AN2CHD U1259 ( .I1(n1657), .I2(n1656), .O(n1658) );
  ND2CHD U1260 ( .I1(n1852), .I2(rkey_next[23]), .O(n1657) );
  ND2CHD U1261 ( .I1(n1807), .I2(Kin[23]), .O(n1656) );
  ND2CHD U1262 ( .I1(n1347), .I2(n1605), .O(n466) );
  AN2CHD U1263 ( .I1(n1346), .I2(n1345), .O(n1347) );
  ND2CHD U1264 ( .I1(rkey_next[23]), .I2(n1584), .O(n1345) );
  ND2CHD U1265 ( .I1(n1852), .I2(rkey_next[39]), .O(n1346) );
  AN2CHD U1266 ( .I1(n1650), .I2(n1649), .O(n1651) );
  AN2CHD U1267 ( .I1(n1645), .I2(n1644), .O(n1646) );
  AN2CHD U1268 ( .I1(n1641), .I2(n1640), .O(n1642) );
  ND2CHD U1269 ( .I1(n1852), .I2(rkey_next[26]), .O(n1641) );
  ND2CHD U1270 ( .I1(n1807), .I2(Kin[26]), .O(n1640) );
  ND2CHD U1271 ( .I1(n1516), .I2(n1599), .O(n470) );
  AN2CHD U1272 ( .I1(n1515), .I2(n1514), .O(n1516) );
  ND2CHD U1273 ( .I1(rkey_next[26]), .I2(n1584), .O(n1514) );
  ND2CHD U1274 ( .I1(n1852), .I2(rkey_next[42]), .O(n1515) );
  AN2CHD U1275 ( .I1(n1634), .I2(n1633), .O(n1635) );
  ND2CHD U1276 ( .I1(n1851), .I2(key[45]), .O(n1634) );
  AN2CHD U1277 ( .I1(n1625), .I2(n1624), .O(n1626) );
  ND2CHD U1278 ( .I1(n1852), .I2(rkey_next[29]), .O(n1625) );
  ND2CHD U1279 ( .I1(n1540), .I2(n1593), .O(n474) );
  AN2CHD U1280 ( .I1(n1539), .I2(n1538), .O(n1540) );
  ND2CHD U1281 ( .I1(rkey_next[29]), .I2(n1584), .O(n1538) );
  ND2CHD U1282 ( .I1(n1852), .I2(rkey_next[45]), .O(n1539) );
  ND2CHD U1283 ( .I1(n1510), .I2(n1509), .O(n476) );
  ND2CHD U1284 ( .I1(n1852), .I2(rkey_next[16]), .O(n1510) );
  ND2CHD U1285 ( .I1(n1546), .I2(n1619), .O(n477) );
  AN2CHD U1286 ( .I1(n1545), .I2(n1544), .O(n1546) );
  ND2CHD U1287 ( .I1(rkey_next[16]), .I2(n1584), .O(n1544) );
  ND2CHD U1288 ( .I1(n1852), .I2(rkey_next[32]), .O(n1545) );
  AN2CHD U1289 ( .I1(n1549), .I2(n1587), .O(n1550) );
  ND2CHD U1290 ( .I1(rkey_next[32]), .I2(n1584), .O(n1549) );
  INVDHD U1291 ( .I(n869), .O(n824) );
  OR2EHD U1292 ( .I1(n764), .I2(n766), .O(n620) );
  AN2CHD U1293 ( .I1(n942), .I2(n941), .O(n623) );
  INVDHD U1294 ( .I(n797), .O(n1164) );
  ND2DHD U1295 ( .I1(n800), .I2(n799), .O(n797) );
  AN2CHD U1296 ( .I1(n1110), .I2(n782), .O(n624) );
  INVKHD U1297 ( .I(n631), .O(n718) );
  AN2HHD U1298 ( .I1(n819), .I2(n946), .O(n820) );
  INVGHD U1299 ( .I(n792), .O(n1156) );
  XNR3EHD U1300 ( .I1(n1242), .I2(n627), .I3(n1099), .O(n1128) );
  XNR3EHD U1301 ( .I1(n929), .I2(n928), .I3(n962), .O(n930) );
  OA22EHD U1302 ( .A1(n1285), .A2(n699), .B1(n1287), .B2(\keyexpantion/N26 ), 
        .O(n1286) );
  XNR2KHD U1303 ( .I1(n1174), .I2(n1173), .O(n699) );
  OAI12CHD U1304 ( .B1(n1226), .B2(n1225), .A1(n628), .O(n629) );
  INVGHD U1305 ( .I(n1276), .O(n628) );
  XOR2HHD U1306 ( .I1(n956), .I2(n927), .O(n772) );
  XOR2HHD U1307 ( .I1(n1110), .I2(n636), .O(n927) );
  NR2GHD U1308 ( .I1(n869), .I2(n822), .O(n819) );
  INVGHD U1309 ( .I(n1058), .O(n709) );
  XNR2KHD U1310 ( .I1(n615), .I2(n629), .O(n677) );
  ND2KHD U1311 ( .I1(n630), .I2(n682), .O(n721) );
  ND3EHD U1312 ( .I1(n814), .I2(n812), .I3(n813), .O(n630) );
  INVGHD U1313 ( .I(n1057), .O(n708) );
  INVGHD U1314 ( .I(n1109), .O(n666) );
  INVHHD U1315 ( .I(n1287), .O(n631) );
  ND2KHD U1316 ( .I1(n1168), .I2(n1169), .O(n1183) );
  AN2HHD U1317 ( .I1(n840), .I2(n820), .O(n841) );
  INVLHD U1318 ( .I(n1329), .O(n935) );
  XNR3EHD U1319 ( .I1(n1021), .I2(n1029), .I3(n1031), .O(n1058) );
  NR2GHD U1320 ( .I1(n791), .I2(n808), .O(n807) );
  INVCKGHD U1321 ( .I(n1219), .O(n1220) );
  XNR2HHD U1322 ( .I1(n1189), .I2(n1199), .O(n1197) );
  INVDHD U1323 ( .I(n1291), .O(n725) );
  OAI22CHD U1324 ( .A1(n1060), .A2(n633), .B1(n644), .B2(n1054), .O(n1086) );
  ND3EHD U1325 ( .I1(n648), .I2(n647), .I3(n646), .O(n633) );
  XOR2HHD U1326 ( .I1(n1060), .I2(n633), .O(n643) );
  INVGHD U1327 ( .I(n634), .O(n1229) );
  ND2HHD U1328 ( .I1(n635), .I2(n1177), .O(n634) );
  ND2HHD U1329 ( .I1(n635), .I2(n752), .O(n684) );
  ND2HHD U1330 ( .I1(n1176), .I2(n635), .O(n1184) );
  ND2KHD U1331 ( .I1(n1170), .I2(n1171), .O(n635) );
  XNR2HHD U1332 ( .I1(n957), .I2(n959), .O(n956) );
  XOR2HHD U1333 ( .I1(n952), .I2(n1143), .O(n636) );
  XOR2HHD U1334 ( .I1(n1563), .I2(n773), .O(n1143) );
  ND2HHD U1335 ( .I1(n640), .I2(n639), .O(n1287) );
  ND3EHD U1336 ( .I1(n658), .I2(n1183), .I3(n1184), .O(n639) );
  ND2HHD U1337 ( .I1(n642), .I2(n641), .O(n640) );
  INVDHD U1338 ( .I(n1184), .O(n641) );
  ND2HHD U1339 ( .I1(n721), .I2(n1177), .O(n658) );
  ND2HHD U1340 ( .I1(n643), .I2(n722), .O(n776) );
  OAI22CHD U1341 ( .A1(n1086), .A2(n1085), .B1(n722), .B2(n643), .O(n707) );
  ND2DHD U1342 ( .I1(n1086), .I2(n1085), .O(n809) );
  MAOI1CHD U1343 ( .A1(n1052), .A2(n645), .B1(n1040), .B2(n1047), .O(n644) );
  ND3CHD U1344 ( .I1(n1053), .I2(n1078), .I3(n1054), .O(n646) );
  ND3EHD U1345 ( .I1(n645), .I2(n1052), .I3(n1051), .O(n647) );
  ND2DHD U1346 ( .I1(n697), .I2(n696), .O(n648) );
  XNR2HHD U1347 ( .I1(n1041), .I2(n649), .O(n1060) );
  XOR2HHD U1348 ( .I1(n1042), .I2(n1043), .O(n649) );
  XOR2HHD U1349 ( .I1(n626), .I2(n1547), .O(n1296) );
  ND2HHD U1350 ( .I1(n654), .I2(n650), .O(n1547) );
  ND3EHD U1351 ( .I1(n653), .I2(n652), .I3(n651), .O(n650) );
  ND2HHD U1352 ( .I1(n729), .I2(n1293), .O(n651) );
  ND2HHD U1353 ( .I1(n731), .I2(n730), .O(n653) );
  ND2HHD U1354 ( .I1(n656), .I2(n655), .O(n654) );
  NR2GHD U1355 ( .I1(n726), .I2(n723), .O(n655) );
  OAI12CHD U1356 ( .B1(n732), .B2(n677), .A1(n676), .O(n656) );
  ND2HHD U1357 ( .I1(n1059), .I2(n657), .O(n705) );
  XOR2HHD U1358 ( .I1(n1159), .I2(n1160), .O(n657) );
  NR2BHD U1359 ( .I1(n1175), .I2(n658), .O(n1182) );
  ND2HHD U1360 ( .I1(n1040), .I2(n1047), .O(n1052) );
  OA12HHD U1361 ( .B1(n661), .B2(n660), .A1(n659), .O(n1040) );
  ND2HHD U1362 ( .I1(n1089), .I2(n704), .O(n659) );
  NR2GHD U1363 ( .I1(n1045), .I2(n1089), .O(n661) );
  OAI12CHD U1364 ( .B1(n1056), .B2(n1055), .A1(n815), .O(n1057) );
  XOR2HHD U1365 ( .I1(n1020), .I2(n662), .O(n1055) );
  XOR2HHD U1366 ( .I1(n1016), .I2(n1017), .O(n662) );
  XOR2HHD U1367 ( .I1(n1093), .I2(n1010), .O(n1016) );
  ND2HHD U1368 ( .I1(n664), .I2(n663), .O(n1003) );
  ND3EHD U1369 ( .I1(n622), .I2(n1002), .I3(n999), .O(n663) );
  ND2HHD U1370 ( .I1(n747), .I2(n1041), .O(n664) );
  NR2IHD U1371 ( .I1(n618), .I2(n667), .O(n1157) );
  XOR2HHD U1372 ( .I1(n1167), .I2(n668), .O(n1169) );
  ND2KHD U1373 ( .I1(n692), .I2(n688), .O(n668) );
  MUX2HHD U1374 ( .A(n672), .B(n671), .S(n996), .O(n669) );
  ND2HHD U1375 ( .I1(n985), .I2(n670), .O(n996) );
  ND3CHD U1376 ( .I1(n974), .I2(n973), .I3(rnd[16]), .O(n670) );
  XOR2HHD U1377 ( .I1(n976), .I2(n1319), .O(n985) );
  ND2HHD U1378 ( .I1(n1136), .I2(n993), .O(n672) );
  MXL2CHD U1379 ( .A(n674), .B(n675), .S(n1136), .OB(n673) );
  INVLHD U1380 ( .I(n994), .O(n1136) );
  XNR2HHD U1381 ( .I1(n972), .I2(n971), .O(n994) );
  NR2CHD U1382 ( .I1(n675), .I2(n993), .O(n674) );
  INVCKGHD U1383 ( .I(n995), .O(n675) );
  INVCKIHD U1384 ( .I(n677), .O(n1283) );
  ND2DHD U1385 ( .I1(n1228), .I2(n677), .O(n676) );
  ND2HHD U1386 ( .I1(n677), .I2(n1286), .O(n730) );
  ND2HHD U1387 ( .I1(n679), .I2(n678), .O(n1202) );
  AO12CHD U1388 ( .B1(n974), .B2(n824), .A1(n1350), .O(n679) );
  ND2HHD U1389 ( .I1(n680), .I2(n1291), .O(n1282) );
  INVCKIHD U1390 ( .I(n1288), .O(n680) );
  AN2HHD U1391 ( .I1(n1285), .I2(\keyexpantion/N26 ), .O(n1288) );
  XNR2CHD U1392 ( .I1(n1254), .I2(n1115), .O(n1253) );
  XNR2HHD U1393 ( .I1(n1115), .I2(n1118), .O(n1163) );
  ND2HHD U1394 ( .I1(n1225), .I2(n683), .O(n1173) );
  ND2HHD U1395 ( .I1(n721), .I2(n1229), .O(n1225) );
  NR2GHD U1396 ( .I1(n811), .I2(n807), .O(n682) );
  ND2HHD U1397 ( .I1(n684), .I2(n1176), .O(n1222) );
  ND2HHD U1398 ( .I1(n695), .I2(n1172), .O(n1176) );
  ND2HHD U1399 ( .I1(n685), .I2(n1553), .O(n803) );
  ND2HHD U1400 ( .I1(n806), .I2(n805), .O(n685) );
  ND2HHD U1401 ( .I1(n686), .I2(n797), .O(n805) );
  ND2HHD U1402 ( .I1(n1160), .I2(n687), .O(n806) );
  ND2HHD U1403 ( .I1(n756), .I2(n759), .O(n1160) );
  MUX2HHD U1404 ( .A(n690), .B(n689), .S(n785), .O(n688) );
  OAI12CHD U1405 ( .B1(n1022), .B2(n893), .A1(n894), .O(n689) );
  ND2CHD U1406 ( .I1(n1022), .I2(n893), .O(n691) );
  MUX2HHD U1407 ( .A(n693), .B(n617), .S(n1024), .O(n692) );
  ND2CHD U1408 ( .I1(n785), .I2(n1022), .O(n693) );
  XNR2KHD U1409 ( .I1(n1138), .I2(n825), .O(n785) );
  XOR2HHD U1410 ( .I1(n720), .I2(n694), .O(n1073) );
  ND2HHD U1411 ( .I1(n974), .I2(n839), .O(n694) );
  INVGHD U1412 ( .I(n1170), .O(n695) );
  XOR2HHD U1413 ( .I1(n1158), .I2(n1157), .O(n1170) );
  ND2DHD U1414 ( .I1(n1051), .I2(n1053), .O(n696) );
  NR2GHD U1415 ( .I1(n988), .I2(n1000), .O(n1043) );
  ND2HHD U1416 ( .I1(n1001), .I2(n998), .O(n1042) );
  INVMHD U1417 ( .I(n699), .O(n1291) );
  OA22EHD U1418 ( .A1(n1227), .A2(n699), .B1(n1287), .B2(n1857), .O(n1228) );
  INVCHD U1419 ( .I(n1072), .O(n703) );
  INVGHD U1420 ( .I(n1089), .O(n1077) );
  INVCHD U1421 ( .I(n1090), .O(n704) );
  NR2EHD U1422 ( .I1(n707), .I2(n791), .O(n814) );
  ND2HHD U1423 ( .I1(n706), .I2(n705), .O(n791) );
  ND2HHD U1424 ( .I1(n709), .I2(n708), .O(n706) );
  XOR2HHD U1425 ( .I1(n1055), .I2(n1056), .O(n1085) );
  AN2HHD U1426 ( .I1(n741), .I2(n619), .O(n1059) );
  ND3EHD U1427 ( .I1(n714), .I2(n713), .I3(n710), .O(n734) );
  MXL2CHD U1428 ( .A(n1271), .B(n1275), .S(n1274), .OB(n713) );
  MAOI1CHD U1429 ( .A1(n1274), .A2(n1273), .B1(n1278), .B2(n1277), .O(n714) );
  INVCHD U1430 ( .I(n1234), .O(n1248) );
  OAI22CHD U1431 ( .A1(n1265), .A2(n1264), .B1(n715), .B2(n1263), .O(n1266) );
  XNR2HHD U1432 ( .I1(n717), .I2(n716), .O(n1264) );
  XNR2HHD U1433 ( .I1(n1249), .I2(n1234), .O(n716) );
  INVDHD U1434 ( .I(n1263), .O(n717) );
  AN2HHD U1435 ( .I1(n1287), .I2(\keyexpantion/N26 ), .O(n728) );
  XOR2EHD U1436 ( .I1(n1036), .I2(n1037), .O(n720) );
  NR2EHD U1437 ( .I1(rnd[4]), .I2(rnd[3]), .O(n969) );
  ND3CHD U1438 ( .I1(n721), .I2(n1272), .I3(n1230), .O(n1231) );
  XNR2HHD U1439 ( .I1(n1185), .I2(n721), .O(n1285) );
  NR2BHD U1440 ( .I1(n721), .I2(n1179), .O(n1180) );
  ND2HHD U1441 ( .I1(n736), .I2(n1084), .O(n722) );
  ND2HHD U1442 ( .I1(n725), .I2(n1279), .O(n724) );
  ND2HHD U1443 ( .I1(n734), .I2(n727), .O(n726) );
  ND3EHD U1444 ( .I1(n728), .I2(n1291), .I3(n1280), .O(n727) );
  ND2HHD U1445 ( .I1(n1290), .I2(n1289), .O(n729) );
  ND2HHD U1446 ( .I1(n1284), .I2(n1283), .O(n731) );
  OAI22CHD U1447 ( .A1(n1291), .A2(n1187), .B1(n1186), .B2(n718), .O(n732) );
  OAI12CHD U1448 ( .B1(n614), .B2(n798), .A1(n733), .O(n760) );
  XOR2HHD U1449 ( .I1(n1252), .I2(n1026), .O(n1021) );
  XOR2HHD U1450 ( .I1(n1095), .I2(n1114), .O(n1026) );
  XOR2HHD U1451 ( .I1(n1561), .I2(n794), .O(n1114) );
  ND2HHD U1452 ( .I1(n1214), .I2(n1190), .O(n1095) );
  INVCHD U1453 ( .I(n1280), .O(n735) );
  ND2DHD U1454 ( .I1(n1087), .I2(n1088), .O(n736) );
  XNR3EHD U1455 ( .I1(n1080), .I2(n1079), .I3(n1078), .O(n1088) );
  XOR2HHD U1456 ( .I1(n909), .I2(n737), .O(n771) );
  XOR2CHD U1457 ( .I1(n737), .I2(n870), .O(n897) );
  ND2HHD U1458 ( .I1(n974), .I2(n973), .O(n737) );
  ND2DHD U1459 ( .I1(n738), .I2(n1042), .O(n747) );
  INVGHD U1460 ( .I(n1043), .O(n738) );
  XOR2HHD U1461 ( .I1(n986), .I2(n771), .O(n1062) );
  ND2HHD U1462 ( .I1(n743), .I2(n742), .O(n1102) );
  ND2HHD U1463 ( .I1(n1119), .I2(n1096), .O(n743) );
  ND2HHD U1464 ( .I1(n744), .I2(n1211), .O(n1119) );
  ND2HHD U1465 ( .I1(n1144), .I2(rnd[28]), .O(n744) );
  ND2CHD U1466 ( .I1(n968), .I2(n969), .O(n746) );
  INVCKGHD U1467 ( .I(n1183), .O(n752) );
  ND2HHD U1468 ( .I1(n803), .I2(n804), .O(n1168) );
  XNR3EHD U1469 ( .I1(n922), .I2(n921), .I3(n772), .O(n1158) );
  XNR2HHD U1470 ( .I1(n1027), .I2(n753), .O(n1161) );
  ND2HHD U1471 ( .I1(n1009), .I2(n1008), .O(n753) );
  ND2HHD U1472 ( .I1(n1291), .I2(n1292), .O(n1293) );
  ND2HHD U1473 ( .I1(n718), .I2(n1281), .O(n1292) );
  NR2GHD U1474 ( .I1(\keyexpantion/N26 ), .I2(n1285), .O(n1281) );
  XOR2HHD U1475 ( .I1(n1122), .I2(n1123), .O(n1126) );
  ND2DHD U1476 ( .I1(n1091), .I2(n755), .O(n1011) );
  ND2DHD U1477 ( .I1(n1093), .I2(n755), .O(n1094) );
  OAI12CHD U1478 ( .B1(n757), .B2(n798), .A1(n797), .O(n756) );
  ND2HHD U1479 ( .I1(n760), .I2(n1164), .O(n759) );
  ND2KHD U1480 ( .I1(n937), .I2(n796), .O(n869) );
  NR2IHD U1481 ( .I1(rnd[11]), .I2(rnd[10]), .O(n796) );
  NR2IHD U1482 ( .I1(rnd[13]), .I2(rnd[12]), .O(n937) );
  ND2HHD U1483 ( .I1(n766), .I2(n765), .O(n1091) );
  ND2HHD U1484 ( .I1(n1010), .I2(n1093), .O(n1012) );
  ND3EHD U1485 ( .I1(n620), .I2(n763), .I3(n761), .O(n1010) );
  ND2DHD U1486 ( .I1(n762), .I2(n982), .O(n761) );
  INVGHD U1487 ( .I(n982), .O(n764) );
  ND3EHD U1488 ( .I1(n940), .I2(n942), .I3(n625), .O(n765) );
  AO12HHD U1489 ( .B1(n623), .B2(n940), .A1(n767), .O(n766) );
  XOR2HHD U1490 ( .I1(n1107), .I2(n1108), .O(n1093) );
  ND2CHD U1491 ( .I1(n946), .I2(n945), .O(n1107) );
  ND2HHD U1492 ( .I1(n768), .I2(n864), .O(n801) );
  ND2HHD U1493 ( .I1(n768), .I2(n908), .O(n783) );
  XOR2HHD U1494 ( .I1(n1188), .I2(n1193), .O(n964) );
  XNR2HHD U1495 ( .I1(n1195), .I2(n769), .O(n1193) );
  XNR3EHD U1496 ( .I1(n1204), .I2(n1198), .I3(n770), .O(n769) );
  XOR2EHD U1497 ( .I1(n1190), .I2(n1205), .O(n770) );
  MAO222CHD U1498 ( .A1(n772), .B1(n962), .C1(n963), .O(n1188) );
  ND2HHD U1499 ( .I1(n1177), .I2(n1183), .O(n1185) );
  OR3HHD U1500 ( .I1(n779), .I2(n778), .I3(n792), .O(n812) );
  ND2HHD U1501 ( .I1(n776), .I2(n777), .O(n792) );
  ND2HHD U1502 ( .I1(n1152), .I2(n1151), .O(n777) );
  NR2CHD U1503 ( .I1(n1150), .I2(n1149), .O(n778) );
  XNR2HHD U1504 ( .I1(n1128), .I2(n1127), .O(n1150) );
  OAI22CHD U1505 ( .A1(n784), .A2(n624), .B1(n781), .B2(n1133), .O(n1122) );
  INVCHD U1506 ( .I(n1132), .O(n781) );
  ND2CHD U1507 ( .I1(n1111), .I2(n1109), .O(n782) );
  XNR2KHD U1508 ( .I1(rnd[27]), .I2(n783), .O(n1110) );
  OAI22CHD U1509 ( .A1(n1112), .A2(n1132), .B1(n1111), .B2(n793), .O(n784) );
  XOR2HHD U1510 ( .I1(n914), .I2(n632), .O(n977) );
  INVGHD U1511 ( .I(n1054), .O(n1051) );
  XNR2KHD U1512 ( .I1(n1032), .I2(n1110), .O(n1054) );
  XOR2HHD U1513 ( .I1(n1130), .I2(n1135), .O(n1032) );
  XOR2HHD U1514 ( .I1(n1557), .I2(n916), .O(n1135) );
  XOR2HHD U1515 ( .I1(n793), .I2(n920), .O(n1130) );
  INVCHD U1516 ( .I(rnd[17]), .O(n793) );
  XOR2HHD U1517 ( .I1(n795), .I2(n1107), .O(n1214) );
  INVCHD U1518 ( .I(rnd[13]), .O(n795) );
  AN2CHD U1519 ( .I1(n796), .I2(n1557), .O(n945) );
  ND2HHD U1520 ( .I1(n917), .I2(n796), .O(n1315) );
  ND2CHD U1521 ( .I1(n946), .I2(n796), .O(n916) );
  XNR3EHD U1522 ( .I1(n1105), .I2(n1092), .I3(n970), .O(n1020) );
  ND2DHD U1523 ( .I1(n1066), .I2(n1025), .O(n799) );
  ND2DHD U1524 ( .I1(n1026), .I2(n1252), .O(n800) );
  XNR2KHD U1525 ( .I1(rnd[30]), .I2(n801), .O(n1250) );
  NR2GHD U1526 ( .I1(n802), .I2(n910), .O(n840) );
  ND2HHD U1527 ( .I1(n936), .I2(n934), .O(n910) );
  NR2EHD U1528 ( .I1(rnd[21]), .I2(rnd[20]), .O(n936) );
  NR2EHD U1529 ( .I1(rnd[23]), .I2(rnd[22]), .O(n872) );
  ND3EHD U1530 ( .I1(n806), .I2(\keyexpantion/N27 ), .I3(n805), .O(n804) );
  ND2KHD U1531 ( .I1(n842), .I2(n933), .O(n975) );
  NR2IHD U1532 ( .I1(rnd[5]), .I2(rnd[4]), .O(n933) );
  NR2IHD U1533 ( .I1(rnd[3]), .I2(rnd[2]), .O(n842) );
  XNR3EHD U1534 ( .I1(n1035), .I2(n990), .I3(n1140), .O(n1078) );
  AN2HHD U1535 ( .I1(n810), .I2(n809), .O(n808) );
  ND2HHD U1536 ( .I1(n1155), .I2(n1156), .O(n813) );
  NR2EHD U1537 ( .I1(n1232), .I2(n1231), .O(n1273) );
  ND2CHD U1538 ( .I1(dat_next[8]), .I2(dat_next[15]), .O(n817) );
  XOR2CHD U1539 ( .I1(dat_next[14]), .I2(Dout[0]), .O(n816) );
  XNR2CHD U1540 ( .I1(n817), .I2(n816), .O(n818) );
  ND2KHD U1541 ( .I1(n840), .I2(n871), .O(n1033) );
  NR2IHD U1542 ( .I1(rnd[9]), .I2(rnd[8]), .O(n1306) );
  NR2IHD U1543 ( .I1(rnd[7]), .I2(rnd[6]), .O(n943) );
  NR2IHD U1544 ( .I1(n932), .I2(n975), .O(n946) );
  INVKHD U1545 ( .I(rnd[15]), .O(n1559) );
  ND2KHD U1546 ( .I1(n1559), .I2(n1350), .O(n868) );
  ND2HHD U1547 ( .I1(n917), .I2(n1305), .O(n822) );
  INVGHD U1548 ( .I(n989), .O(n1138) );
  BUFNHD U1549 ( .I(n946), .O(n974) );
  XNR2KHD U1550 ( .I1(n1556), .I2(n974), .O(n1137) );
  ND2HHD U1551 ( .I1(n1137), .I2(n1038), .O(n912) );
  XOR2HHD U1552 ( .I1(n912), .I2(n1140), .O(n825) );
  INVDHD U1553 ( .I(n1038), .O(n827) );
  XNR2KHD U1554 ( .I1(n827), .I2(n826), .O(n1251) );
  NR2IHD U1555 ( .I1(n878), .I2(n869), .O(n834) );
  ND2DHD U1556 ( .I1(n917), .I2(n1560), .O(n830) );
  ND3CHD U1557 ( .I1(n834), .I2(n832), .I3(n829), .O(n838) );
  ND3CHD U1558 ( .I1(n832), .I2(n943), .I3(n831), .O(n833) );
  INVGHD U1559 ( .I(n834), .O(n835) );
  AN3HHD U1560 ( .I1(n838), .I2(n837), .I3(n836), .O(n1044) );
  INVGHD U1561 ( .I(n1044), .O(n890) );
  XNR2HHD U1562 ( .I1(n890), .I2(n1039), .O(n1244) );
  XNR2KHD U1563 ( .I1(n1251), .I2(n1244), .O(n1022) );
  XNR2KHD U1564 ( .I1(n1564), .I2(n841), .O(n1115) );
  ND3CHD U1565 ( .I1(n935), .I2(n853), .I3(n968), .O(n844) );
  XOR2HHD U1566 ( .I1(n935), .I2(rnd[9]), .O(n845) );
  XOR2EHD U1567 ( .I1(n846), .I2(n845), .O(n1069) );
  INVCHD U1568 ( .I(n1069), .O(n847) );
  ND2DHD U1569 ( .I1(n848), .I2(n847), .O(n850) );
  ND2HHD U1570 ( .I1(n850), .I2(n849), .O(n1024) );
  ND3CHD U1571 ( .I1(n872), .I2(n851), .I3(n1564), .O(n852) );
  XOR2HHD U1572 ( .I1(rnd[4]), .I2(n935), .O(n1215) );
  BUFGHD U1573 ( .I(n933), .O(n915) );
  XOR2CHD U1574 ( .I1(rnd[9]), .I2(rnd[25]), .O(n855) );
  OAI12CHD U1575 ( .B1(n879), .B2(n854), .A1(n855), .O(n859) );
  INVCHD U1576 ( .I(n855), .O(n857) );
  ND3CHD U1577 ( .I1(n857), .I2(n856), .I3(n915), .O(n858) );
  ND3CHD U1578 ( .I1(n859), .I2(n1215), .I3(n858), .O(n860) );
  XOR2HHD U1579 ( .I1(n877), .I2(n862), .O(n883) );
  NR2EHD U1580 ( .I1(rnd[26]), .I2(rnd[27]), .O(n1013) );
  NR2BHD U1581 ( .I1(rnd[28]), .I2(rnd[29]), .O(n863) );
  NR2EHD U1582 ( .I1(n874), .I2(n1033), .O(n864) );
  XOR2HHD U1583 ( .I1(n883), .I2(n1250), .O(n1023) );
  INVDHD U1584 ( .I(n1023), .O(n894) );
  NR2BHD U1585 ( .I1(rnd[10]), .I2(rnd[7]), .O(n865) );
  ND3CHD U1586 ( .I1(n872), .I2(n871), .I3(n1568), .O(n873) );
  OR3CHD U1587 ( .I1(n874), .I2(n910), .I3(n873), .O(n875) );
  NR2EHD U1588 ( .I1(n879), .I2(n878), .O(n880) );
  XNR2EHD U1589 ( .I1(n1555), .I2(n880), .O(n1240) );
  ND2HHD U1590 ( .I1(n1240), .I2(n1215), .O(n1071) );
  INVCHD U1591 ( .I(n1071), .O(n881) );
  INVDHD U1592 ( .I(n883), .O(n884) );
  INVDHD U1593 ( .I(n890), .O(n1045) );
  MAO222CHD U1594 ( .A1(n1022), .B1(n894), .C1(n893), .O(n895) );
  INVCHD U1595 ( .I(n897), .O(n900) );
  NR2EHD U1596 ( .I1(rnd[31]), .I2(n898), .O(n987) );
  INVCHD U1597 ( .I(n987), .O(n899) );
  ND2HHD U1598 ( .I1(n999), .I2(n901), .O(n963) );
  XOR2HHD U1599 ( .I1(rnd[2]), .I2(n963), .O(n922) );
  ND2HHD U1600 ( .I1(n907), .I2(n925), .O(n921) );
  NR2EHD U1601 ( .I1(rnd[26]), .I2(n1033), .O(n908) );
  ND3EHD U1602 ( .I1(n935), .I2(n915), .I3(n914), .O(n971) );
  ND2CHD U1603 ( .I1(n937), .I2(n909), .O(n918) );
  ND2DHD U1604 ( .I1(n946), .I2(n919), .O(n920) );
  XNR3EHD U1605 ( .I1(n950), .I2(n1135), .I3(n666), .O(n957) );
  INVDHD U1606 ( .I(n1158), .O(n931) );
  INVGHD U1607 ( .I(n927), .O(n961) );
  XOR2HHD U1608 ( .I1(n963), .I2(n961), .O(n928) );
  OA22EHD U1609 ( .A1(n1157), .A2(n931), .B1(n930), .B2(rnd[2]), .O(n965) );
  NR2EHD U1610 ( .I1(n932), .I2(n1315), .O(n942) );
  NR2EHD U1611 ( .I1(n1316), .I2(n975), .O(n944) );
  XOR2EHD U1612 ( .I1(n1144), .I2(n1210), .O(n1198) );
  INVCHD U1613 ( .I(n1013), .O(n947) );
  ND2HHD U1614 ( .I1(n955), .I2(n954), .O(n1204) );
  ND2HHD U1615 ( .I1(n967), .I2(n966), .O(n1223) );
  ND2HHD U1616 ( .I1(n1230), .I2(n1223), .O(n1174) );
  ND2HHD U1617 ( .I1(n997), .I2(n1136), .O(n980) );
  ND2HHD U1618 ( .I1(n1143), .I2(n994), .O(n978) );
  ND2HHD U1619 ( .I1(n978), .I2(n1131), .O(n979) );
  ND2HHD U1620 ( .I1(n980), .I2(n979), .O(n1017) );
  INVDHD U1621 ( .I(n1130), .O(n1109) );
  ND2HHD U1622 ( .I1(n1012), .I2(n1011), .O(n1027) );
  XOR2HHD U1623 ( .I1(n614), .I2(n1161), .O(n1031) );
  INVCHD U1624 ( .I(rnd[28]), .O(n1567) );
  ND2CHD U1625 ( .I1(n1013), .I2(n1567), .O(n1014) );
  INVDHD U1626 ( .I(n1016), .O(n1019) );
  INVGHD U1627 ( .I(n1017), .O(n1018) );
  MAO222HHD U1628 ( .A1(n1020), .B1(n1019), .C1(n1018), .O(n1029) );
  XNR3EHD U1629 ( .I1(n1024), .I2(n1023), .I3(n1022), .O(n1159) );
  INVCHD U1630 ( .I(n1095), .O(n1025) );
  XOR2HHD U1631 ( .I1(n1028), .I2(n1029), .O(n1030) );
  OAI12CHD U1632 ( .B1(n1034), .B2(n1033), .A1(n1565), .O(n1035) );
  XNR2KHD U1633 ( .I1(\keyexpantion/N26 ), .I2(n1137), .O(n1089) );
  XOR2CHD U1634 ( .I1(rnd[5]), .I2(rnd[15]), .O(n1036) );
  NR2CHD U1635 ( .I1(n1046), .I2(n1045), .O(n1076) );
  OAI12CHD U1636 ( .B1(n1566), .B2(n1098), .A1(n1074), .O(n1080) );
  OAI12CHD U1637 ( .B1(n1077), .B2(n1076), .A1(n1075), .O(n1079) );
  INVCHD U1638 ( .I(n1082), .O(n1083) );
  ND2DHD U1639 ( .I1(n1081), .I2(n1083), .O(n1084) );
  XOR2HHD U1640 ( .I1(n1088), .I2(n1087), .O(n1152) );
  XNR3EHD U1641 ( .I1(n1090), .I2(n1250), .I3(n1089), .O(n1101) );
  AN2HHD U1642 ( .I1(n1095), .I2(n1094), .O(n1117) );
  NR2BHD U1643 ( .I1(n1117), .I2(n1118), .O(n1097) );
  XOR2HHD U1644 ( .I1(n1101), .I2(n1102), .O(n1127) );
  BUFIHD U1645 ( .I(n1114), .O(n1247) );
  XNR3EHD U1646 ( .I1(n1116), .I2(n1247), .I3(n1115), .O(n1123) );
  XNR3EHD U1647 ( .I1(n1121), .I2(n1120), .I3(n1119), .O(n1129) );
  ND2CHD U1648 ( .I1(n1124), .I2(n1123), .O(n1125) );
  INVCHD U1649 ( .I(n1149), .O(n1154) );
  OAI22CHD U1650 ( .A1(n1154), .A2(n1153), .B1(n1152), .B2(n1151), .O(n1155)
         );
  INVDHD U1651 ( .I(n1171), .O(n1172) );
  MXL2CHD U1652 ( .A(n1177), .B(n1183), .S(n1184), .OB(n1181) );
  INVCHD U1653 ( .I(n1185), .O(n1178) );
  AN2EHD U1654 ( .I1(n1184), .I2(n1178), .O(n1179) );
  OA13EHD U1655 ( .B1(n1182), .B2(n1181), .B3(n1180), .A1(\keyexpantion/N26 ), 
        .O(n1187) );
  INVDHD U1656 ( .I(n1281), .O(n1186) );
  INVCHD U1657 ( .I(n1188), .O(n1194) );
  INVCHD U1658 ( .I(n1198), .O(n1189) );
  XOR2HHD U1659 ( .I1(n1195), .I2(n1197), .O(n1192) );
  INVCHD U1660 ( .I(n1190), .O(n1191) );
  OA22EHD U1661 ( .A1(n1194), .A2(n1193), .B1(n1192), .B2(n1191), .O(n1219) );
  INVDHD U1662 ( .I(n1195), .O(n1196) );
  ND2HHD U1663 ( .I1(n1197), .I2(n1196), .O(n1201) );
  ND2DHD U1664 ( .I1(n1199), .I2(n1198), .O(n1200) );
  XNR2EHD U1665 ( .I1(n1247), .I2(n1245), .O(n1234) );
  ND2DHD U1666 ( .I1(n1205), .I2(n1204), .O(n1209) );
  ND2HHD U1667 ( .I1(n1209), .I2(n1208), .O(n1233) );
  XNR3EHD U1668 ( .I1(n1249), .I2(n1215), .I3(n1263), .O(n1216) );
  XOR2HHD U1669 ( .I1(n1235), .I2(n1236), .O(n1218) );
  ND2HHD U1670 ( .I1(n1219), .I2(n1218), .O(n1272) );
  INVDHD U1671 ( .I(n1218), .O(n1221) );
  ND2DHD U1672 ( .I1(n1221), .I2(n1220), .O(n1270) );
  ND2HHD U1673 ( .I1(n1222), .I2(n1230), .O(n1224) );
  ND2HHD U1674 ( .I1(n1224), .I2(n1223), .O(n1276) );
  INVCHD U1675 ( .I(n1230), .O(n1226) );
  ND2CHD U1676 ( .I1(n1285), .I2(n1857), .O(n1227) );
  INVDHD U1677 ( .I(n1229), .O(n1232) );
  OAI22CHD U1678 ( .A1(n1239), .A2(n1238), .B1(n1237), .B2(n1236), .O(n1269)
         );
  ND2CHD U1679 ( .I1(n1202), .I2(n1240), .O(n1241) );
  XOR2EHD U1680 ( .I1(n1242), .I2(n1241), .O(n1243) );
  OAI22CHD U1681 ( .A1(n1249), .A2(n1248), .B1(n1247), .B2(n1246), .O(n1261)
         );
  OAI22CHD U1682 ( .A1(n1257), .A2(n1256), .B1(n1255), .B2(n1254), .O(n1258)
         );
  XNR2CHD U1683 ( .I1(n1259), .I2(n1258), .O(n1260) );
  XNR2EHD U1684 ( .I1(n1267), .I2(n1266), .O(n1268) );
  XOR2HHD U1685 ( .I1(n1269), .I2(n1268), .O(n1274) );
  INVDHD U1686 ( .I(n1276), .O(n1277) );
  INVGHD U1687 ( .I(n718), .O(n1279) );
  ND2HHD U1688 ( .I1(n1292), .I2(n1282), .O(n1284) );
  ND2DHD U1689 ( .I1(n1288), .I2(n718), .O(n1290) );
  ND2HHD U1690 ( .I1(n1296), .I2(n1572), .O(n1300) );
  ND2HHD U1691 ( .I1(n1300), .I2(n1299), .O(n500) );
  NR2BHD U1692 ( .I1(rnd[31]), .I2(sel), .O(n1302) );
  ND2CHD U1693 ( .I1(n1302), .I2(n1301), .O(n1322) );
  NR2BHD U1694 ( .I1(rnd[28]), .I2(\keyexpantion/N27 ), .O(n1303) );
  ND2CHD U1695 ( .I1(n1304), .I2(n1303), .O(n1321) );
  NR2BHD U1696 ( .I1(n1308), .I2(n1307), .O(n1314) );
  AN4CHD U1697 ( .I1(n1312), .I2(n1311), .I3(n1310), .I4(n1309), .O(n1313) );
  AN2CHD U1698 ( .I1(n1314), .I2(n1313), .O(n1318) );
  ND3CHD U1699 ( .I1(n1319), .I2(n1318), .I3(n1317), .O(n1320) );
  NR3BHD U1700 ( .I1(n1322), .I2(n1321), .I3(n1320), .O(n1323) );
  MAOI1CHD U1701 ( .A1(EN), .A2(n1323), .B1(BSY), .B2(EN), .O(n480) );
  OA22CHD U1702 ( .A1(n1584), .A2(sel), .B1(Dvld), .B2(EN), .O(n481) );
  INVCHD U1703 ( .I(n1573), .O(n1324) );
  ND2CHD U1704 ( .I1(\keyexpantion/N26 ), .I2(n1324), .O(n1326) );
  ND2CHD U1705 ( .I1(rnd[31]), .I2(EN), .O(n1325) );
  AO12CHD U1706 ( .B1(Kvld), .B2(n1584), .A1(n1807), .O(n483) );
  AOI22BHD U1707 ( .A1(Kin[17]), .A2(n1807), .B1(rkey_next[1]), .B2(n1584), 
        .O(n1331) );
  MXL2CHD U1708 ( .A(n1350), .B(n1559), .S(n1570), .OB(n596) );
  AOI22BHD U1709 ( .A1(Din[18]), .A2(n1573), .B1(dat_next[2]), .B2(n1571), .O(
        n1359) );
  INVCHD U1710 ( .I(rkey_next[37]), .O(n1744) );
  INVCHD U1711 ( .I(rkey_next[2]), .O(n1764) );
  AOI22BHD U1712 ( .A1(rkey_next[2]), .A2(rkey_next[37]), .B1(n1744), .B2(
        n1764), .O(n1412) );
  INVCHD U1713 ( .I(n1412), .O(n1352) );
  INVCHD U1714 ( .I(rkey[2]), .O(n1769) );
  INVCHD U1715 ( .I(rkey_next[38]), .O(n1825) );
  INVCHD U1716 ( .I(rkey_next[3]), .O(n1842) );
  AOI22BHD U1717 ( .A1(rkey_next[3]), .A2(rkey_next[38]), .B1(n1825), .B2(
        n1842), .O(n1380) );
  MUX2CHD U1718 ( .A(rkey[2]), .B(n1769), .S(n1380), .O(n1351) );
  XOR2CHD U1719 ( .I1(dat_next[0]), .I2(Dout[2]), .O(n1355) );
  ND2CHD U1720 ( .I1(dat_next[10]), .I2(dat_next[1]), .O(n1354) );
  ND2CHD U1721 ( .I1(n1354), .I2(n1355), .O(n1353) );
  OAI12CHD U1722 ( .B1(n1355), .B2(n1354), .A1(n1353), .O(n1357) );
  ND2CHD U1723 ( .I1(n1758), .I2(n1357), .O(n1356) );
  OAI112BHD U1724 ( .C1(n1758), .C2(n1357), .A1(n1572), .B1(n1356), .O(n1358)
         );
  AOI22BHD U1725 ( .A1(Din[27]), .A2(n1573), .B1(dat_next[11]), .B2(n1571), 
        .O(n1369) );
  INVCHD U1726 ( .I(rkey_next[46]), .O(n1696) );
  INVCHD U1727 ( .I(rkey_next[11]), .O(n1716) );
  AOI22BHD U1728 ( .A1(rkey_next[11]), .A2(rkey_next[46]), .B1(n1696), .B2(
        n1716), .O(n1400) );
  INVCHD U1729 ( .I(n1400), .O(n1361) );
  INVCHD U1730 ( .I(rkey[11]), .O(n1721) );
  INVCHD U1731 ( .I(rkey_next[47]), .O(n1776) );
  INVCHD U1732 ( .I(rkey_next[12]), .O(n1796) );
  AOI22BHD U1733 ( .A1(rkey_next[12]), .A2(rkey_next[47]), .B1(n1776), .B2(
        n1796), .O(n1390) );
  MUX2CHD U1734 ( .A(rkey[11]), .B(n1721), .S(n1390), .O(n1360) );
  INVCHD U1735 ( .I(dat_next[10]), .O(n1365) );
  MAOI1CHD U1736 ( .A1(dat_next[9]), .A2(Dout[11]), .B1(Dout[11]), .B2(
        dat_next[9]), .O(n1364) );
  INVCHD U1737 ( .I(dat_next[3]), .O(n1363) );
  OAI12CHD U1738 ( .B1(n1365), .B2(n1363), .A1(n1364), .O(n1362) );
  OAI13BHD U1739 ( .B1(n1365), .B2(n1364), .B3(n1363), .A1(n1362), .O(n1367)
         );
  ND2CHD U1740 ( .I1(n1710), .I2(n1367), .O(n1366) );
  OAI112BHD U1741 ( .C1(n1710), .C2(n1367), .A1(n1572), .B1(n1366), .O(n1368)
         );
  AOI22BHD U1742 ( .A1(Din[23]), .A2(n1573), .B1(dat_next[7]), .B2(n1571), .O(
        n1378) );
  INVCHD U1743 ( .I(rkey_next[42]), .O(n1639) );
  INVCHD U1744 ( .I(rkey_next[7]), .O(n1659) );
  AOI22BHD U1745 ( .A1(rkey_next[7]), .A2(rkey_next[42]), .B1(n1639), .B2(
        n1659), .O(n1433) );
  INVCHD U1746 ( .I(n1433), .O(n1371) );
  INVCHD U1747 ( .I(rkey[7]), .O(n1664) );
  INVCHD U1748 ( .I(rkey_next[43]), .O(n1712) );
  INVCHD U1749 ( .I(rkey_next[8]), .O(n1732) );
  AOI22BHD U1750 ( .A1(rkey_next[8]), .A2(rkey_next[43]), .B1(n1712), .B2(
        n1732), .O(n1486) );
  MUX2CHD U1751 ( .A(rkey[7]), .B(n1664), .S(n1486), .O(n1370) );
  INVCHD U1752 ( .I(dat_next[15]), .O(n1374) );
  MAOI1CHD U1753 ( .A1(dat_next[5]), .A2(Dout[7]), .B1(Dout[7]), .B2(
        dat_next[5]), .O(n1373) );
  INVCHD U1754 ( .I(dat_next[6]), .O(n1477) );
  OAI12CHD U1755 ( .B1(n1374), .B2(n1477), .A1(n1373), .O(n1372) );
  OAI13BHD U1756 ( .B1(n1374), .B2(n1373), .B3(n1477), .A1(n1372), .O(n1376)
         );
  ND2CHD U1757 ( .I1(n1653), .I2(n1376), .O(n1375) );
  OAI112BHD U1758 ( .C1(n1653), .C2(n1376), .A1(n1572), .B1(n1375), .O(n1377)
         );
  AOI22BHD U1759 ( .A1(Din[19]), .A2(n1573), .B1(dat_next[3]), .B2(n1571), .O(
        n1388) );
  INVCHD U1760 ( .I(n1380), .O(n1381) );
  INVCHD U1761 ( .I(rkey[3]), .O(n1850) );
  INVCHD U1762 ( .I(rkey_next[39]), .O(n1655) );
  INVCHD U1763 ( .I(rkey_next[4]), .O(n1672) );
  AOI22BHD U1764 ( .A1(rkey_next[4]), .A2(rkey_next[39]), .B1(n1655), .B2(
        n1672), .O(n1464) );
  MUX2CHD U1765 ( .A(rkey[3]), .B(n1850), .S(n1464), .O(n1379) );
  MAOI1CHD U1766 ( .A1(dat_next[1]), .A2(Dout[3]), .B1(Dout[3]), .B2(
        dat_next[1]), .O(n1384) );
  ND2CHD U1767 ( .I1(dat_next[11]), .I2(dat_next[2]), .O(n1383) );
  ND2CHD U1768 ( .I1(n1383), .I2(n1384), .O(n1382) );
  OAI12CHD U1769 ( .B1(n1384), .B2(n1383), .A1(n1382), .O(n1386) );
  ND2CHD U1770 ( .I1(n1511), .I2(n1386), .O(n1385) );
  OAI112BHD U1771 ( .C1(n1511), .C2(n1386), .A1(n1572), .B1(n1385), .O(n1387)
         );
  AOI22BHD U1772 ( .A1(Din[28]), .A2(n1573), .B1(dat_next[12]), .B2(n1571), 
        .O(n1399) );
  INVCHD U1773 ( .I(n1390), .O(n1391) );
  INVCHD U1774 ( .I(rkey[12]), .O(n1801) );
  MUX2CHD U1775 ( .A(rkey[12]), .B(n1801), .S(n1453), .O(n1389) );
  INVCHD U1776 ( .I(dat_next[11]), .O(n1395) );
  MAOI1CHD U1777 ( .A1(dat_next[10]), .A2(Dout[12]), .B1(Dout[12]), .B2(
        dat_next[10]), .O(n1394) );
  INVCHD U1778 ( .I(dat_next[4]), .O(n1393) );
  OAI12CHD U1779 ( .B1(n1395), .B2(n1393), .A1(n1394), .O(n1392) );
  OAI13BHD U1780 ( .B1(n1395), .B2(n1394), .B3(n1393), .A1(n1392), .O(n1397)
         );
  ND2CHD U1781 ( .I1(n1790), .I2(n1397), .O(n1396) );
  OAI112BHD U1782 ( .C1(n1790), .C2(n1397), .A1(n1572), .B1(n1396), .O(n1398)
         );
  AOI22BHD U1783 ( .A1(Din[26]), .A2(n1573), .B1(dat_next[10]), .B2(n1571), 
        .O(n1410) );
  INVCHD U1784 ( .I(rkey_next[45]), .O(n1623) );
  INVCHD U1785 ( .I(rkey_next[10]), .O(n1643) );
  AOI22BHD U1786 ( .A1(rkey_next[10]), .A2(rkey_next[45]), .B1(n1623), .B2(
        n1643), .O(n1422) );
  INVCHD U1787 ( .I(n1422), .O(n1402) );
  INVCHD U1788 ( .I(rkey[10]), .O(n1648) );
  MUX2CHD U1789 ( .A(rkey[10]), .B(n1648), .S(n1400), .O(n1401) );
  INVCHD U1790 ( .I(dat_next[9]), .O(n1406) );
  MAOI1CHD U1791 ( .A1(dat_next[8]), .A2(Dout[10]), .B1(Dout[10]), .B2(
        dat_next[8]), .O(n1405) );
  INVCHD U1792 ( .I(dat_next[2]), .O(n1404) );
  OAI12CHD U1793 ( .B1(n1406), .B2(n1404), .A1(n1405), .O(n1403) );
  OAI13BHD U1794 ( .B1(n1406), .B2(n1405), .B3(n1404), .A1(n1403), .O(n1408)
         );
  ND2CHD U1795 ( .I1(n1637), .I2(n1408), .O(n1407) );
  OAI112BHD U1796 ( .C1(n1637), .C2(n1408), .A1(n1572), .B1(n1407), .O(n1409)
         );
  AOI22BHD U1797 ( .A1(Din[17]), .A2(n1573), .B1(dat_next[1]), .B2(n1571), .O(
        n1421) );
  INVCHD U1798 ( .I(n1411), .O(n1414) );
  INVCHD U1799 ( .I(rkey[1]), .O(n1689) );
  MAOI1CHD U1800 ( .A1(dat_next[15]), .A2(Dout[1]), .B1(Dout[1]), .B2(
        dat_next[15]), .O(n1417) );
  ND2CHD U1801 ( .I1(dat_next[0]), .I2(dat_next[9]), .O(n1416) );
  ND2CHD U1802 ( .I1(n1416), .I2(n1417), .O(n1415) );
  OAI12CHD U1803 ( .B1(n1417), .B2(n1416), .A1(n1415), .O(n1419) );
  ND2CHD U1804 ( .I1(n1682), .I2(n1419), .O(n1418) );
  OAI112BHD U1805 ( .C1(n1682), .C2(n1419), .A1(n1572), .B1(n1418), .O(n1420)
         );
  AOI22BHD U1806 ( .A1(Din[25]), .A2(n1573), .B1(dat_next[9]), .B2(n1571), .O(
        n1432) );
  INVCHD U1807 ( .I(rkey_next[44]), .O(n1792) );
  INVCHD U1808 ( .I(rkey_next[9]), .O(n1813) );
  AOI22BHD U1809 ( .A1(rkey_next[9]), .A2(rkey_next[44]), .B1(n1792), .B2(
        n1813), .O(n1484) );
  INVCHD U1810 ( .I(n1484), .O(n1424) );
  INVCHD U1811 ( .I(rkey[9]), .O(n1818) );
  MUX2CHD U1812 ( .A(rkey[9]), .B(n1818), .S(n1422), .O(n1423) );
  INVCHD U1813 ( .I(dat_next[8]), .O(n1428) );
  MAOI1CHD U1814 ( .A1(dat_next[7]), .A2(Dout[9]), .B1(Dout[9]), .B2(
        dat_next[7]), .O(n1427) );
  INVCHD U1815 ( .I(dat_next[1]), .O(n1426) );
  OAI12CHD U1816 ( .B1(n1428), .B2(n1426), .A1(n1427), .O(n1425) );
  OAI13BHD U1817 ( .B1(n1428), .B2(n1427), .B3(n1426), .A1(n1425), .O(n1430)
         );
  ND2CHD U1818 ( .I1(n1806), .I2(n1430), .O(n1429) );
  OAI112BHD U1819 ( .C1(n1806), .C2(n1430), .A1(n1572), .B1(n1429), .O(n1431)
         );
  AOI22BHD U1820 ( .A1(Din[22]), .A2(n1573), .B1(dat_next[6]), .B2(n1571), .O(
        n1441) );
  INVCHD U1821 ( .I(rkey_next[41]), .O(n1809) );
  INVCHD U1822 ( .I(rkey_next[6]), .O(n1829) );
  AOI22BHD U1823 ( .A1(rkey_next[6]), .A2(rkey_next[41]), .B1(n1809), .B2(
        n1829), .O(n1442) );
  INVCHD U1824 ( .I(n1442), .O(n1435) );
  INVCHD U1825 ( .I(rkey[6]), .O(n1834) );
  MUX2CHD U1826 ( .A(rkey[6]), .B(n1834), .S(n1433), .O(n1434) );
  INVCHD U1827 ( .I(dat_next[14]), .O(n1501) );
  MAOI1CHD U1828 ( .A1(dat_next[4]), .A2(Dout[6]), .B1(Dout[6]), .B2(
        dat_next[4]), .O(n1437) );
  INVCHD U1829 ( .I(dat_next[5]), .O(n1455) );
  OAI12CHD U1830 ( .B1(n1501), .B2(n1455), .A1(n1437), .O(n1436) );
  OAI13BHD U1831 ( .B1(n1501), .B2(n1437), .B3(n1455), .A1(n1436), .O(n1439)
         );
  ND2CHD U1832 ( .I1(n1823), .I2(n1439), .O(n1438) );
  OAI112BHD U1833 ( .C1(n1823), .C2(n1439), .A1(n1572), .B1(n1438), .O(n1440)
         );
  AOI22BHD U1834 ( .A1(Din[21]), .A2(n1573), .B1(dat_next[5]), .B2(n1571), .O(
        n1451) );
  INVCHD U1835 ( .I(rkey_next[40]), .O(n1728) );
  INVCHD U1836 ( .I(rkey_next[5]), .O(n1748) );
  AOI22BHD U1837 ( .A1(rkey_next[5]), .A2(rkey_next[40]), .B1(n1728), .B2(
        n1748), .O(n1462) );
  INVCHD U1838 ( .I(n1462), .O(n1444) );
  INVCHD U1839 ( .I(rkey[5]), .O(n1753) );
  MUX2CHD U1840 ( .A(rkey[5]), .B(n1753), .S(n1442), .O(n1443) );
  MAOI1CHD U1841 ( .A1(dat_next[3]), .A2(Dout[5]), .B1(Dout[5]), .B2(
        dat_next[3]), .O(n1447) );
  ND2CHD U1842 ( .I1(dat_next[13]), .I2(dat_next[4]), .O(n1446) );
  ND2CHD U1843 ( .I1(n1446), .I2(n1447), .O(n1445) );
  OAI12CHD U1844 ( .B1(n1447), .B2(n1446), .A1(n1445), .O(n1449) );
  ND2CHD U1845 ( .I1(n1742), .I2(n1449), .O(n1448) );
  OAI112BHD U1846 ( .C1(n1742), .C2(n1449), .A1(n1572), .B1(n1448), .O(n1450)
         );
  AOI22BHD U1847 ( .A1(Din[29]), .A2(n1573), .B1(dat_next[13]), .B2(n1571), 
        .O(n1461) );
  INVCHD U1848 ( .I(rkey[13]), .O(n1632) );
  INVCHD U1849 ( .I(rkey_next[33]), .O(n1684) );
  INVCHD U1850 ( .I(rkey_next[14]), .O(n1700) );
  AOI22BHD U1851 ( .A1(rkey_next[14]), .A2(rkey_next[33]), .B1(n1684), .B2(
        n1700), .O(n1474) );
  INVCHD U1852 ( .I(dat_next[12]), .O(n1457) );
  MAOI1CHD U1853 ( .A1(dat_next[11]), .A2(Dout[13]), .B1(Dout[13]), .B2(
        dat_next[11]), .O(n1456) );
  OAI12CHD U1854 ( .B1(n1457), .B2(n1455), .A1(n1456), .O(n1454) );
  OAI13BHD U1855 ( .B1(n1457), .B2(n1456), .B3(n1455), .A1(n1454), .O(n1459)
         );
  ND2CHD U1856 ( .I1(n1621), .I2(n1459), .O(n1458) );
  OAI112BHD U1857 ( .C1(n1621), .C2(n1459), .A1(n1572), .B1(n1458), .O(n1460)
         );
  AOI22BHD U1858 ( .A1(Din[20]), .A2(n1573), .B1(dat_next[4]), .B2(n1571), .O(
        n1472) );
  INVCHD U1859 ( .I(n1464), .O(n1465) );
  INVCHD U1860 ( .I(rkey[4]), .O(n1677) );
  MUX2CHD U1861 ( .A(rkey[4]), .B(n1677), .S(n1462), .O(n1463) );
  MAOI1CHD U1862 ( .A1(dat_next[2]), .A2(Dout[4]), .B1(Dout[4]), .B2(
        dat_next[2]), .O(n1468) );
  ND2CHD U1863 ( .I1(dat_next[12]), .I2(dat_next[3]), .O(n1467) );
  ND2CHD U1864 ( .I1(n1467), .I2(n1468), .O(n1466) );
  OAI12CHD U1865 ( .B1(n1468), .B2(n1467), .A1(n1466), .O(n1470) );
  ND2CHD U1866 ( .I1(n1506), .I2(n1470), .O(n1469) );
  OAI112BHD U1867 ( .C1(n1506), .C2(n1470), .A1(n1572), .B1(n1469), .O(n1471)
         );
  AOI22BHD U1868 ( .A1(dat_next[14]), .A2(n1571), .B1(n1573), .B2(Din[30]), 
        .O(n1483) );
  INVCHD U1869 ( .I(n1474), .O(n1475) );
  INVCHD U1870 ( .I(rkey[14]), .O(n1705) );
  INVCHD U1871 ( .I(rkey_next[34]), .O(n1760) );
  INVCHD U1872 ( .I(rkey_next[15]), .O(n1780) );
  AOI22BHD U1873 ( .A1(rkey_next[15]), .A2(rkey_next[34]), .B1(n1760), .B2(
        n1780), .O(n1495) );
  MUX2CHD U1874 ( .A(rkey[14]), .B(n1705), .S(n1495), .O(n1473) );
  INVCHD U1875 ( .I(dat_next[13]), .O(n1479) );
  MAOI1CHD U1876 ( .A1(dat_next[12]), .A2(Dout[14]), .B1(Dout[14]), .B2(
        dat_next[12]), .O(n1478) );
  OAI12CHD U1877 ( .B1(n1479), .B2(n1477), .A1(n1478), .O(n1476) );
  OAI13BHD U1878 ( .B1(n1479), .B2(n1478), .B3(n1477), .A1(n1476), .O(n1481)
         );
  ND2CHD U1879 ( .I1(n1694), .I2(n1481), .O(n1480) );
  OAI112BHD U1880 ( .C1(n1694), .C2(n1481), .A1(n1572), .B1(n1480), .O(n1482)
         );
  AOI22BHD U1881 ( .A1(dat_next[8]), .A2(n1571), .B1(n1573), .B2(Din[24]), .O(
        n1494) );
  INVCHD U1882 ( .I(n1486), .O(n1487) );
  INVCHD U1883 ( .I(rkey[8]), .O(n1737) );
  MUX2CHD U1884 ( .A(rkey[8]), .B(n1737), .S(n1484), .O(n1485) );
  MAOI1CHD U1885 ( .A1(dat_next[6]), .A2(Dout[8]), .B1(Dout[8]), .B2(
        dat_next[6]), .O(n1490) );
  INVCHD U1886 ( .I(dat_next[0]), .O(n1488) );
  INVCHD U1887 ( .I(dat_next[7]), .O(n1499) );
  OR2CHD U1888 ( .I1(n1488), .I2(n1499), .O(n1489) );
  XNR2CHD U1889 ( .I1(n1490), .I2(n1489), .O(n1492) );
  ND2CHD U1890 ( .I1(n1726), .I2(n1492), .O(n1491) );
  OAI112BHD U1891 ( .C1(n1726), .C2(n1492), .A1(n1572), .B1(n1491), .O(n1493)
         );
  AOI22BHD U1892 ( .A1(dat_next[15]), .A2(n1571), .B1(n1573), .B2(Din[31]), 
        .O(n1505) );
  MAOI1CHD U1893 ( .A1(n1495), .A2(rkey[15]), .B1(rkey[15]), .B2(n1495), .O(
        n1496) );
  MAOI1CHD U1894 ( .A1(dat_next[13]), .A2(Dout[15]), .B1(Dout[15]), .B2(
        dat_next[13]), .O(n1500) );
  OAI12CHD U1895 ( .B1(n1501), .B2(n1499), .A1(n1500), .O(n1498) );
  OAI13BHD U1896 ( .B1(n1501), .B2(n1500), .B3(n1499), .A1(n1498), .O(n1503)
         );
  ND2CHD U1897 ( .I1(n1774), .I2(n1503), .O(n1502) );
  OAI112BHD U1898 ( .C1(n1774), .C2(n1503), .A1(n1572), .B1(n1502), .O(n1504)
         );
  AOI22BHD U1899 ( .A1(Kin[52]), .A2(n1807), .B1(rkey_next[36]), .B2(n1584), 
        .O(n1507) );
  AOI22BHD U1900 ( .A1(Kin[16]), .A2(n1807), .B1(rkey_next[0]), .B2(n1584), 
        .O(n1509) );
  AOI22BHD U1901 ( .A1(Kin[51]), .A2(n1807), .B1(rkey_next[35]), .B2(n1584), 
        .O(n1512) );
  XNR2HHD U1902 ( .I1(n1548), .I2(n1547), .O(n1552) );
  OAI12CHD U1903 ( .B1(n1552), .B2(n1551), .A1(n1550), .O(n478) );
  MXL2CHD U1904 ( .A(n1857), .B(n1553), .S(n1570), .OB(n610) );
  MXL2CHD U1905 ( .A(n1553), .B(n1579), .S(n1570), .OB(n609) );
  MXL2CHD U1906 ( .A(n1554), .B(n1555), .S(n1570), .OB(n602) );
  MXL2CHD U1907 ( .A(n1555), .B(n1556), .S(n1570), .OB(n601) );
  MXL2CHD U1908 ( .A(n1556), .B(n1558), .S(n1570), .OB(n600) );
  MXL2CHD U1909 ( .A(n1558), .B(n1557), .S(n1570), .OB(n599) );
  MXL2CHD U1910 ( .A(n1559), .B(n909), .S(n1570), .OB(n595) );
  MXL2CHD U1911 ( .A(n788), .B(n1563), .S(n1570), .OB(n589) );
  MXL2CHD U1912 ( .A(n1564), .B(n1566), .S(n1570), .OB(n586) );
  MXL2CHD U1913 ( .A(n1566), .B(n1565), .S(n1570), .OB(n585) );
  MXL2CHD U1914 ( .A(n1567), .B(n1569), .S(n1570), .OB(n582) );
  MXL2CHD U1915 ( .A(n1569), .B(n1568), .S(n1570), .OB(n581) );
  MUX2CHD U1916 ( .A(sel), .B(rnd[31]), .S(EN), .O(n482) );
  ND2CHD U1917 ( .I1(n1573), .I2(Din[0]), .O(n1574) );
  ND3CHD U1918 ( .I1(n1576), .I2(n1575), .I3(n1574), .O(n516) );
  INVCHD U1919 ( .I(rkey_next[0]), .O(n1582) );
  AOI22BHD U1920 ( .A1(n1845), .A2(key[48]), .B1(n1851), .B2(key[32]), .O(
        n1581) );
  AOI22BHD U1921 ( .A1(n1807), .A2(Kin[0]), .B1(rkey[0]), .B2(n1584), .O(n1580) );
  OAI112BHD U1922 ( .C1(n1551), .C2(n1582), .A1(n1581), .B1(n1580), .O(n1586)
         );
  NR3BHD U1923 ( .I1(Krdy), .I2(n1857), .I3(n1584), .O(n1843) );
  AOI22BHD U1924 ( .A1(n1844), .A2(key[16]), .B1(n1843), .B2(key[0]), .O(n1585) );
  OR2B1CHD U1925 ( .I1(n1586), .B1(n1585), .O(n479) );
  INVCHD U1926 ( .I(key[48]), .O(n1588) );
  OAI12CHD U1927 ( .B1(n1807), .B2(n1588), .A1(n1587), .O(n565) );
  INVCHD U1928 ( .I(key[47]), .O(n1590) );
  OAI12CHD U1929 ( .B1(n1807), .B2(n1590), .A1(n1589), .O(n564) );
  INVCHD U1930 ( .I(key[46]), .O(n1592) );
  OAI12CHD U1931 ( .B1(n1807), .B2(n1592), .A1(n1591), .O(n563) );
  INVCHD U1932 ( .I(key[45]), .O(n1594) );
  OAI12CHD U1933 ( .B1(n1807), .B2(n1594), .A1(n1593), .O(n562) );
  INVCHD U1934 ( .I(key[44]), .O(n1596) );
  OAI12CHD U1935 ( .B1(n1807), .B2(n1596), .A1(n1595), .O(n561) );
  INVCHD U1936 ( .I(key[43]), .O(n1598) );
  OAI12CHD U1937 ( .B1(n1807), .B2(n1598), .A1(n1597), .O(n560) );
  INVCHD U1938 ( .I(key[42]), .O(n1600) );
  OAI12CHD U1939 ( .B1(n1807), .B2(n1600), .A1(n1599), .O(n559) );
  INVCHD U1940 ( .I(key[41]), .O(n1602) );
  OAI12CHD U1941 ( .B1(n1807), .B2(n1602), .A1(n1601), .O(n558) );
  INVCHD U1942 ( .I(key[40]), .O(n1604) );
  OAI12CHD U1943 ( .B1(n1807), .B2(n1604), .A1(n1603), .O(n557) );
  INVCHD U1944 ( .I(key[39]), .O(n1606) );
  OAI12CHD U1945 ( .B1(n1807), .B2(n1606), .A1(n1605), .O(n556) );
  INVCHD U1946 ( .I(key[38]), .O(n1608) );
  OAI12CHD U1947 ( .B1(n1807), .B2(n1608), .A1(n1607), .O(n555) );
  INVCHD U1948 ( .I(key[37]), .O(n1610) );
  OAI12CHD U1949 ( .B1(n1807), .B2(n1610), .A1(n1609), .O(n554) );
  INVCHD U1950 ( .I(key[36]), .O(n1612) );
  OAI12CHD U1951 ( .B1(n1807), .B2(n1612), .A1(n1611), .O(n553) );
  INVCHD U1952 ( .I(key[35]), .O(n1614) );
  OAI12CHD U1953 ( .B1(n1807), .B2(n1614), .A1(n1613), .O(n552) );
  INVCHD U1954 ( .I(key[34]), .O(n1616) );
  OAI12CHD U1955 ( .B1(n1807), .B2(n1616), .A1(n1615), .O(n551) );
  INVCHD U1956 ( .I(key[33]), .O(n1618) );
  OAI12CHD U1957 ( .B1(n1807), .B2(n1618), .A1(n1617), .O(n550) );
  INVCHD U1958 ( .I(key[32]), .O(n1620) );
  OAI12CHD U1959 ( .B1(n1807), .B2(n1620), .A1(n1619), .O(n549) );
  AOI22BHD U1960 ( .A1(n1807), .A2(Kin[61]), .B1(n1621), .B2(n1852), .O(n1622)
         );
  OAI12CHD U1961 ( .B1(EN), .B2(n1623), .A1(n1622), .O(n475) );
  INVCHD U1962 ( .I(rkey_next[13]), .O(n1627) );
  OAI12CHD U1963 ( .B1(EN), .B2(n1627), .A1(n1626), .O(n473) );
  AOI22BHD U1964 ( .A1(n1844), .A2(key[29]), .B1(n1843), .B2(key[13]), .O(
        n1631) );
  OAI112BHD U1965 ( .C1(EN), .C2(n1632), .A1(n1631), .B1(n1630), .O(n1636) );
  OR2B1CHD U1966 ( .I1(n1636), .B1(n1635), .O(n472) );
  AOI22BHD U1967 ( .A1(n1807), .A2(Kin[58]), .B1(n1637), .B2(n1852), .O(n1638)
         );
  OAI12CHD U1968 ( .B1(EN), .B2(n1639), .A1(n1638), .O(n471) );
  OAI12CHD U1969 ( .B1(EN), .B2(n1643), .A1(n1642), .O(n469) );
  AOI22BHD U1970 ( .A1(n1844), .A2(key[26]), .B1(n1843), .B2(key[10]), .O(
        n1647) );
  ND2CHD U1971 ( .I1(n1807), .I2(Kin[10]), .O(n1644) );
  OAI112BHD U1972 ( .C1(EN), .C2(n1648), .A1(n1647), .B1(n1646), .O(n1652) );
  OR2B1CHD U1973 ( .I1(n1652), .B1(n1651), .O(n468) );
  AOI22BHD U1974 ( .A1(n1807), .A2(Kin[55]), .B1(n1653), .B2(n1852), .O(n1654)
         );
  OAI12CHD U1975 ( .B1(EN), .B2(n1655), .A1(n1654), .O(n467) );
  OAI12CHD U1976 ( .B1(EN), .B2(n1659), .A1(n1658), .O(n465) );
  AOI22BHD U1977 ( .A1(n1844), .A2(key[23]), .B1(n1843), .B2(key[7]), .O(n1663) );
  OAI112BHD U1978 ( .C1(EN), .C2(n1664), .A1(n1663), .B1(n1662), .O(n1668) );
  OR2B1CHD U1979 ( .I1(n1668), .B1(n1667), .O(n464) );
  OAI12CHD U1980 ( .B1(EN), .B2(n1672), .A1(n1671), .O(n461) );
  AOI22BHD U1981 ( .A1(n1844), .A2(key[20]), .B1(n1843), .B2(key[4]), .O(n1676) );
  ND2CHD U1982 ( .I1(n1807), .I2(Kin[4]), .O(n1673) );
  OAI112BHD U1983 ( .C1(EN), .C2(n1677), .A1(n1676), .B1(n1675), .O(n1681) );
  OR2B1CHD U1984 ( .I1(n1681), .B1(n1680), .O(n460) );
  AOI22BHD U1985 ( .A1(n1807), .A2(Kin[49]), .B1(n1682), .B2(n1852), .O(n1683)
         );
  OAI12CHD U1986 ( .B1(EN), .B2(n1684), .A1(n1683), .O(n459) );
  AOI22BHD U1987 ( .A1(n1844), .A2(key[17]), .B1(n1843), .B2(key[1]), .O(n1688) );
  ND2CHD U1988 ( .I1(n1807), .I2(Kin[1]), .O(n1685) );
  OAI112BHD U1989 ( .C1(EN), .C2(n1689), .A1(n1688), .B1(n1687), .O(n1693) );
  OR2B1CHD U1990 ( .I1(n1693), .B1(n1692), .O(n456) );
  AOI22BHD U1991 ( .A1(n1807), .A2(Kin[62]), .B1(n1694), .B2(n1852), .O(n1695)
         );
  OAI12CHD U1992 ( .B1(EN), .B2(n1696), .A1(n1695), .O(n455) );
  OAI12CHD U1993 ( .B1(EN), .B2(n1700), .A1(n1699), .O(n453) );
  AOI22BHD U1994 ( .A1(n1844), .A2(key[30]), .B1(n1843), .B2(key[14]), .O(
        n1704) );
  ND2CHD U1995 ( .I1(n1807), .I2(Kin[14]), .O(n1701) );
  OAI112BHD U1996 ( .C1(EN), .C2(n1705), .A1(n1704), .B1(n1703), .O(n1709) );
  OR2B1CHD U1997 ( .I1(n1709), .B1(n1708), .O(n452) );
  AOI22BHD U1998 ( .A1(n1807), .A2(Kin[59]), .B1(n1710), .B2(n1852), .O(n1711)
         );
  OAI12CHD U1999 ( .B1(EN), .B2(n1712), .A1(n1711), .O(n451) );
  OAI12CHD U2000 ( .B1(EN), .B2(n1716), .A1(n1715), .O(n449) );
  AOI22BHD U2001 ( .A1(n1844), .A2(key[27]), .B1(n1843), .B2(key[11]), .O(
        n1720) );
  ND2CHD U2002 ( .I1(n1807), .I2(Kin[11]), .O(n1717) );
  OAI112BHD U2003 ( .C1(EN), .C2(n1721), .A1(n1720), .B1(n1719), .O(n1725) );
  OR2B1CHD U2004 ( .I1(n1725), .B1(n1724), .O(n448) );
  AOI22BHD U2005 ( .A1(n1807), .A2(Kin[56]), .B1(n1726), .B2(n1852), .O(n1727)
         );
  OAI12CHD U2006 ( .B1(EN), .B2(n1728), .A1(n1727), .O(n447) );
  OAI12CHD U2007 ( .B1(EN), .B2(n1732), .A1(n1731), .O(n445) );
  AOI22BHD U2008 ( .A1(n1844), .A2(key[24]), .B1(n1843), .B2(key[8]), .O(n1736) );
  OAI112BHD U2009 ( .C1(EN), .C2(n1737), .A1(n1736), .B1(n1735), .O(n1741) );
  OR2B1CHD U2010 ( .I1(n1741), .B1(n1740), .O(n444) );
  AOI22BHD U2011 ( .A1(n1807), .A2(Kin[53]), .B1(n1742), .B2(n1852), .O(n1743)
         );
  OAI12CHD U2012 ( .B1(EN), .B2(n1744), .A1(n1743), .O(n443) );
  OAI12CHD U2013 ( .B1(EN), .B2(n1748), .A1(n1747), .O(n441) );
  AOI22BHD U2014 ( .A1(n1844), .A2(key[21]), .B1(n1843), .B2(key[5]), .O(n1752) );
  ND2CHD U2015 ( .I1(n1807), .I2(Kin[5]), .O(n1749) );
  OAI112BHD U2016 ( .C1(EN), .C2(n1753), .A1(n1752), .B1(n1751), .O(n1757) );
  OR2B1CHD U2017 ( .I1(n1757), .B1(n1756), .O(n440) );
  AOI22BHD U2018 ( .A1(n1807), .A2(Kin[50]), .B1(n1758), .B2(n1852), .O(n1759)
         );
  OAI12CHD U2019 ( .B1(EN), .B2(n1760), .A1(n1759), .O(n439) );
  OAI12CHD U2020 ( .B1(EN), .B2(n1764), .A1(n1763), .O(n437) );
  AOI22BHD U2021 ( .A1(n1844), .A2(key[18]), .B1(n1843), .B2(key[2]), .O(n1768) );
  OAI112BHD U2022 ( .C1(EN), .C2(n1769), .A1(n1768), .B1(n1767), .O(n1773) );
  OR2B1CHD U2023 ( .I1(n1773), .B1(n1772), .O(n436) );
  AOI22BHD U2024 ( .A1(n1807), .A2(Kin[63]), .B1(n1774), .B2(n1852), .O(n1775)
         );
  OAI12CHD U2025 ( .B1(EN), .B2(n1776), .A1(n1775), .O(n435) );
  OAI12CHD U2026 ( .B1(EN), .B2(n1780), .A1(n1779), .O(n433) );
  INVCHD U2027 ( .I(rkey[15]), .O(n1785) );
  AOI22BHD U2028 ( .A1(n1844), .A2(key[31]), .B1(n1843), .B2(key[15]), .O(
        n1784) );
  OAI112BHD U2029 ( .C1(EN), .C2(n1785), .A1(n1784), .B1(n1783), .O(n1789) );
  OR2B1CHD U2030 ( .I1(n1789), .B1(n1788), .O(n432) );
  AOI22BHD U2031 ( .A1(n1807), .A2(Kin[60]), .B1(n1790), .B2(n1852), .O(n1791)
         );
  OAI12CHD U2032 ( .B1(EN), .B2(n1792), .A1(n1791), .O(n431) );
  OAI12CHD U2033 ( .B1(EN), .B2(n1796), .A1(n1795), .O(n429) );
  AOI22BHD U2034 ( .A1(n1844), .A2(key[28]), .B1(n1843), .B2(key[12]), .O(
        n1800) );
  OAI112BHD U2035 ( .C1(EN), .C2(n1801), .A1(n1800), .B1(n1799), .O(n1805) );
  OR2B1CHD U2036 ( .I1(n1805), .B1(n1804), .O(n428) );
  AOI22BHD U2037 ( .A1(n1807), .A2(Kin[57]), .B1(n1806), .B2(n1852), .O(n1808)
         );
  OAI12CHD U2038 ( .B1(EN), .B2(n1809), .A1(n1808), .O(n427) );
  OAI12CHD U2039 ( .B1(EN), .B2(n1813), .A1(n1812), .O(n425) );
  AOI22BHD U2040 ( .A1(n1844), .A2(key[25]), .B1(n1843), .B2(key[9]), .O(n1817) );
  ND2CHD U2041 ( .I1(n1807), .I2(Kin[9]), .O(n1814) );
  OAI112BHD U2042 ( .C1(EN), .C2(n1818), .A1(n1817), .B1(n1816), .O(n1822) );
  OR2B1CHD U2043 ( .I1(n1822), .B1(n1821), .O(n424) );
  AOI22BHD U2044 ( .A1(n1807), .A2(Kin[54]), .B1(n1823), .B2(n1852), .O(n1824)
         );
  OAI12CHD U2045 ( .B1(EN), .B2(n1825), .A1(n1824), .O(n423) );
  OAI12CHD U2046 ( .B1(EN), .B2(n1829), .A1(n1828), .O(n421) );
  AOI22BHD U2047 ( .A1(n1844), .A2(key[22]), .B1(n1843), .B2(key[6]), .O(n1833) );
  ND2CHD U2048 ( .I1(n1807), .I2(Kin[6]), .O(n1830) );
  OAI112BHD U2049 ( .C1(EN), .C2(n1834), .A1(n1833), .B1(n1832), .O(n1838) );
  OR2B1CHD U2050 ( .I1(n1838), .B1(n1837), .O(n420) );
  OAI12CHD U2051 ( .B1(EN), .B2(n1842), .A1(n1841), .O(n417) );
  AOI22BHD U2052 ( .A1(n1844), .A2(key[19]), .B1(n1843), .B2(key[3]), .O(n1849) );
  OAI112BHD U2053 ( .C1(EN), .C2(n1850), .A1(n1849), .B1(n1848), .O(n1856) );
  OR2B1CHD U2054 ( .I1(n1856), .B1(n1855), .O(n416) );
endmodule

